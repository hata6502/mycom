iconv input.asm -f utf8 -t sjis > input.c
gcc -E -P input.c > input_pre.asm
rm input.c
./asm < input_pre.asm
is_word(IS_ADD, 3), 	-- 256
is_word(IS_ADD, 3), 	-- 257
is_word(IS_ADD, 3), 	-- 258
is_word(IS_ADD, 3), 	-- 259
is_word(IS_ADD, 3), 	-- 260
is_word(IS_ADD, 3), 	-- 261
is_word(IS_ADD, 3), 	-- 262
is_word(IS_ADD, 3), 	-- 263
is_word(IS_ADD, 3), 	-- 264
is_word(IS_ADD, 3), 	-- 265
is_word(IS_ADD, 3), 	-- 266
is_word(IS_ADD, 3), 	-- 267
is_word(IS_ADD, 3), 	-- 268
is_word(IS_ADD, 3), 	-- 269
is_word(IS_ADD, 3), 	-- 270
is_word(IS_ADD, 3), 	-- 271
is_word(IS_ADD, 3), 	-- 272
is_word(IS_ADD, 3), 	-- 273
is_word(IS_ADD, 3), 	-- 274
is_word(IS_ADD, 3), 	-- 275
is_word(IS_ADD, 3), 	-- 276
is_word(IS_ADD, 3), 	-- 277
is_word(IS_ADD, 3), 	-- 278
is_word(IS_ADD, 3), 	-- 279
is_word(IS_ADD, 3), 	-- 280
is_word(IS_ADD, 3), 	-- 281
is_word(IS_ADD, 3), 	-- 282
is_word(IS_ADD, 3), 	-- 283
is_word(IS_ADD, 3), 	-- 284
is_word(IS_ADD, 3), 	-- 285
is_word(IS_ADD, 3), 	-- 286
is_word(IS_ADD, 3), 	-- 287
is_word(IS_READ, 767), 	-- 288
is_word(IS_WRITE, 766), 	-- 289
is_word(IS_READ, 765), 	-- 290
is_word(IS_WRITE, 764), 	-- 291
is_word(IS_READ, 763), 	-- 292
is_word(IS_WRITE, 762), 	-- 293
is_word(IS_READ, 761), 	-- 294
is_word(IS_WRITE, 760), 	-- 295
is_word(IS_READ, 11), 	-- 296
is_word(IS_AND, 759), 	-- 297
is_word(IS_BRANCH, 758), 	-- 298
is_word(IS_READ, 757), 	-- 299
is_word(IS_WRITE, 756), 	-- 300
is_word(IS_READ, 755), 	-- 301
is_word(IS_WRITE, 754), 	-- 302
is_word(IS_READ, 11), 	-- 303
is_word(IS_AND, 753), 	-- 304
is_word(IS_BRANCH, 752), 	-- 305
is_word(IS_READ, 751), 	-- 306
is_word(IS_WRITE, 750), 	-- 307
is_word(IS_READ, 749), 	-- 308
is_word(IS_WRITE, 748), 	-- 309
is_word(IS_READ, 11), 	-- 310
is_word(IS_AND, 747), 	-- 311
is_word(IS_BRANCH, 746), 	-- 312
is_word(IS_READ, 9), 	-- 313
is_word(IS_WRITE, 128), 	-- 314
is_word(IS_READ, 128), 	-- 315
is_word(IS_ADD, 745), 	-- 316
is_word(IS_WRITE, 744), 	-- 317
is_word(IS_READ, 743), 	-- 318
is_word(IS_WRITE, 742), 	-- 319
0, 	-- 320
0, 	-- 321
0, 	-- 322
0, 	-- 323
0, 	-- 324
0, 	-- 325
0, 	-- 326
0, 	-- 327
0, 	-- 328
0, 	-- 329
0, 	-- 330
0, 	-- 331
0, 	-- 332
0, 	-- 333
0, 	-- 334
0, 	-- 335
0, 	-- 336
0, 	-- 337
0, 	-- 338
0, 	-- 339
0, 	-- 340
0, 	-- 341
0, 	-- 342
0, 	-- 343
0, 	-- 344
0, 	-- 345
0, 	-- 346
0, 	-- 347
0, 	-- 348
0, 	-- 349
0, 	-- 350
0, 	-- 351
0, 	-- 352
0, 	-- 353
0, 	-- 354
0, 	-- 355
0, 	-- 356
0, 	-- 357
0, 	-- 358
0, 	-- 359
0, 	-- 360
0, 	-- 361
0, 	-- 362
0, 	-- 363
0, 	-- 364
0, 	-- 365
0, 	-- 366
0, 	-- 367
0, 	-- 368
0, 	-- 369
0, 	-- 370
0, 	-- 371
0, 	-- 372
0, 	-- 373
0, 	-- 374
0, 	-- 375
0, 	-- 376
0, 	-- 377
0, 	-- 378
0, 	-- 379
0, 	-- 380
0, 	-- 381
0, 	-- 382
0, 	-- 383
0, 	-- 384
0, 	-- 385
0, 	-- 386
0, 	-- 387
0, 	-- 388
0, 	-- 389
0, 	-- 390
0, 	-- 391
0, 	-- 392
0, 	-- 393
0, 	-- 394
0, 	-- 395
0, 	-- 396
0, 	-- 397
0, 	-- 398
0, 	-- 399
0, 	-- 400
0, 	-- 401
0, 	-- 402
0, 	-- 403
0, 	-- 404
0, 	-- 405
0, 	-- 406
0, 	-- 407
0, 	-- 408
0, 	-- 409
0, 	-- 410
0, 	-- 411
0, 	-- 412
0, 	-- 413
0, 	-- 414
0, 	-- 415
0, 	-- 416
0, 	-- 417
0, 	-- 418
0, 	-- 419
0, 	-- 420
0, 	-- 421
0, 	-- 422
0, 	-- 423
0, 	-- 424
0, 	-- 425
0, 	-- 426
0, 	-- 427
0, 	-- 428
0, 	-- 429
0, 	-- 430
0, 	-- 431
0, 	-- 432
0, 	-- 433
0, 	-- 434
0, 	-- 435
0, 	-- 436
0, 	-- 437
0, 	-- 438
0, 	-- 439
0, 	-- 440
0, 	-- 441
0, 	-- 442
0, 	-- 443
0, 	-- 444
0, 	-- 445
0, 	-- 446
0, 	-- 447
0, 	-- 448
0, 	-- 449
0, 	-- 450
0, 	-- 451
0, 	-- 452
0, 	-- 453
0, 	-- 454
0, 	-- 455
0, 	-- 456
0, 	-- 457
0, 	-- 458
0, 	-- 459
0, 	-- 460
0, 	-- 461
0, 	-- 462
0, 	-- 463
0, 	-- 464
0, 	-- 465
0, 	-- 466
0, 	-- 467
0, 	-- 468
0, 	-- 469
0, 	-- 470
0, 	-- 471
0, 	-- 472
0, 	-- 473
0, 	-- 474
0, 	-- 475
0, 	-- 476
0, 	-- 477
0, 	-- 478
0, 	-- 479
0, 	-- 480
0, 	-- 481
0, 	-- 482
0, 	-- 483
0, 	-- 484
0, 	-- 485
0, 	-- 486
0, 	-- 487
0, 	-- 488
0, 	-- 489
0, 	-- 490
0, 	-- 491
0, 	-- 492
0, 	-- 493
0, 	-- 494
0, 	-- 495
0, 	-- 496
0, 	-- 497
0, 	-- 498
0, 	-- 499
0, 	-- 500
0, 	-- 501
0, 	-- 502
0, 	-- 503
0, 	-- 504
0, 	-- 505
0, 	-- 506
0, 	-- 507
0, 	-- 508
0, 	-- 509
0, 	-- 510
0, 	-- 511
0, 	-- 512
0, 	-- 513
0, 	-- 514
0, 	-- 515
0, 	-- 516
0, 	-- 517
0, 	-- 518
0, 	-- 519
0, 	-- 520
0, 	-- 521
0, 	-- 522
0, 	-- 523
0, 	-- 524
0, 	-- 525
0, 	-- 526
0, 	-- 527
0, 	-- 528
0, 	-- 529
0, 	-- 530
0, 	-- 531
0, 	-- 532
0, 	-- 533
0, 	-- 534
0, 	-- 535
0, 	-- 536
0, 	-- 537
0, 	-- 538
0, 	-- 539
0, 	-- 540
0, 	-- 541
0, 	-- 542
0, 	-- 543
0, 	-- 544
0, 	-- 545
0, 	-- 546
0, 	-- 547
0, 	-- 548
0, 	-- 549
0, 	-- 550
0, 	-- 551
0, 	-- 552
0, 	-- 553
0, 	-- 554
0, 	-- 555
0, 	-- 556
0, 	-- 557
0, 	-- 558
0, 	-- 559
0, 	-- 560
0, 	-- 561
0, 	-- 562
0, 	-- 563
0, 	-- 564
0, 	-- 565
0, 	-- 566
0, 	-- 567
0, 	-- 568
0, 	-- 569
0, 	-- 570
0, 	-- 571
0, 	-- 572
0, 	-- 573
0, 	-- 574
0, 	-- 575
0, 	-- 576
0, 	-- 577
0, 	-- 578
0, 	-- 579
0, 	-- 580
0, 	-- 581
0, 	-- 582
0, 	-- 583
0, 	-- 584
0, 	-- 585
0, 	-- 586
0, 	-- 587
0, 	-- 588
0, 	-- 589
0, 	-- 590
0, 	-- 591
0, 	-- 592
0, 	-- 593
0, 	-- 594
0, 	-- 595
0, 	-- 596
0, 	-- 597
0, 	-- 598
0, 	-- 599
0, 	-- 600
0, 	-- 601
0, 	-- 602
0, 	-- 603
0, 	-- 604
0, 	-- 605
0, 	-- 606
0, 	-- 607
0, 	-- 608
0, 	-- 609
0, 	-- 610
0, 	-- 611
0, 	-- 612
0, 	-- 613
0, 	-- 614
0, 	-- 615
0, 	-- 616
0, 	-- 617
0, 	-- 618
0, 	-- 619
0, 	-- 620
0, 	-- 621
0, 	-- 622
0, 	-- 623
0, 	-- 624
0, 	-- 625
0, 	-- 626
0, 	-- 627
0, 	-- 628
0, 	-- 629
0, 	-- 630
0, 	-- 631
0, 	-- 632
0, 	-- 633
0, 	-- 634
0, 	-- 635
0, 	-- 636
0, 	-- 637
0, 	-- 638
0, 	-- 639
0, 	-- 640
0, 	-- 641
0, 	-- 642
0, 	-- 643
0, 	-- 644
0, 	-- 645
0, 	-- 646
0, 	-- 647
0, 	-- 648
0, 	-- 649
0, 	-- 650
0, 	-- 651
0, 	-- 652
0, 	-- 653
0, 	-- 654
0, 	-- 655
0, 	-- 656
0, 	-- 657
0, 	-- 658
0, 	-- 659
0, 	-- 660
0, 	-- 661
0, 	-- 662
0, 	-- 663
0, 	-- 664
0, 	-- 665
0, 	-- 666
0, 	-- 667
0, 	-- 668
0, 	-- 669
0, 	-- 670
0, 	-- 671
0, 	-- 672
0, 	-- 673
0, 	-- 674
0, 	-- 675
0, 	-- 676
0, 	-- 677
0, 	-- 678
0, 	-- 679
0, 	-- 680
0, 	-- 681
0, 	-- 682
0, 	-- 683
0, 	-- 684
0, 	-- 685
0, 	-- 686
0, 	-- 687
0, 	-- 688
0, 	-- 689
0, 	-- 690
0, 	-- 691
0, 	-- 692
0, 	-- 693
0, 	-- 694
0, 	-- 695
0, 	-- 696
0, 	-- 697
0, 	-- 698
0, 	-- 699
0, 	-- 700
0, 	-- 701
0, 	-- 702
0, 	-- 703
0, 	-- 704
0, 	-- 705
0, 	-- 706
0, 	-- 707
0, 	-- 708
0, 	-- 709
0, 	-- 710
0, 	-- 711
0, 	-- 712
0, 	-- 713
0, 	-- 714
0, 	-- 715
0, 	-- 716
0, 	-- 717
0, 	-- 718
0, 	-- 719
0, 	-- 720
0, 	-- 721
0, 	-- 722
0, 	-- 723
0, 	-- 724
0, 	-- 725
0, 	-- 726
0, 	-- 727
0, 	-- 728
0, 	-- 729
0, 	-- 730
0, 	-- 731
0, 	-- 732
0, 	-- 733
0, 	-- 734
0, 	-- 735
0, 	-- 736
0, 	-- 737
0, 	-- 738
0, 	-- 739
0, 	-- 740
0, 	-- 741
0, 	-- 742
308, 	-- 743
128, 	-- 744
1, 	-- 745
310, 	-- 746
4, 	-- 747
11, 	-- 748
3, 	-- 749
128, 	-- 750
1024, 	-- 751
303, 	-- 752
4, 	-- 753
11, 	-- 754
1, 	-- 755
10, 	-- 756
0, 	-- 757
296, 	-- 758
4, 	-- 759
11, 	-- 760
1, 	-- 761
10, 	-- 762
0, 	-- 763
8, 	-- 764
80, 	-- 765
0, 	-- 766
290	-- 767
