iconv input.asm -f utf8 -t sjis > input.c
gcc -E -P input.c > input_pre.asm
rm input.c
./asm < input_pre.asm
is_word(IS_ADD, 3), 	-- 256
is_word(IS_ADD, 3), 	-- 257
is_word(IS_ADD, 3), 	-- 258
is_word(IS_ADD, 3), 	-- 259
is_word(IS_ADD, 3), 	-- 260
is_word(IS_ADD, 3), 	-- 261
is_word(IS_ADD, 3), 	-- 262
is_word(IS_ADD, 3), 	-- 263
is_word(IS_ADD, 3), 	-- 264
is_word(IS_ADD, 3), 	-- 265
is_word(IS_ADD, 3), 	-- 266
is_word(IS_ADD, 3), 	-- 267
is_word(IS_ADD, 3), 	-- 268
is_word(IS_ADD, 3), 	-- 269
is_word(IS_ADD, 3), 	-- 270
is_word(IS_ADD, 3), 	-- 271
is_word(IS_ADD, 3), 	-- 272
is_word(IS_ADD, 3), 	-- 273
is_word(IS_ADD, 3), 	-- 274
is_word(IS_ADD, 3), 	-- 275
is_word(IS_ADD, 3), 	-- 276
is_word(IS_ADD, 3), 	-- 277
is_word(IS_ADD, 3), 	-- 278
is_word(IS_ADD, 3), 	-- 279
is_word(IS_ADD, 3), 	-- 280
is_word(IS_ADD, 3), 	-- 281
is_word(IS_ADD, 3), 	-- 282
is_word(IS_ADD, 3), 	-- 283
is_word(IS_ADD, 3), 	-- 284
is_word(IS_ADD, 3), 	-- 285
is_word(IS_ADD, 3), 	-- 286
is_word(IS_ADD, 3), 	-- 287
is_word(IS_READ, 767), 	-- 288
is_word(IS_WRITE, 766), 	-- 289
is_word(IS_READ, 66), 	-- 290
is_word(IS_READ, 108), 	-- 291
is_word(IS_READ, 117), 	-- 292
is_word(IS_READ, 101), 	-- 293
is_word(IS_READ, 72), 	-- 294
is_word(IS_READ, 111), 	-- 295
is_word(IS_READ, 111), 	-- 296
is_word(IS_READ, 100), 	-- 297
is_word(IS_READ, 32), 	-- 298
is_word(IS_READ, 67), 	-- 299
is_word(IS_READ, 111), 	-- 300
is_word(IS_READ, 109), 	-- 301
is_word(IS_READ, 112), 	-- 302
is_word(IS_READ, 117), 	-- 303
is_word(IS_READ, 116), 	-- 304
is_word(IS_READ, 101), 	-- 305
is_word(IS_READ, 114), 	-- 306
is_word(IS_READ, 32), 	-- 307
is_word(IS_READ, 32), 	-- 308
is_word(IS_READ, 210), 	-- 309
is_word(IS_READ, 178), 	-- 310
is_word(IS_READ, 219), 	-- 311
is_word(IS_READ, 32), 	-- 312
is_word(IS_READ, 190), 	-- 313
is_word(IS_READ, 178), 	-- 314
is_word(IS_READ, 190), 	-- 315
is_word(IS_READ, 178), 	-- 316
is_word(IS_READ, 32), 	-- 317
is_word(IS_READ, 204), 	-- 318
is_word(IS_READ, 223), 	-- 319
is_word(IS_READ, 219), 	-- 320
is_word(IS_READ, 184), 	-- 321
is_word(IS_READ, 222), 	-- 322
is_word(IS_READ, 215), 	-- 323
is_word(IS_READ, 209), 	-- 324
is_word(IS_READ, 0), 	-- 325
is_word(IS_READ, 219), 	-- 326
is_word(IS_READ, 0), 	-- 327
is_word(IS_READ, 765), 	-- 328
is_word(IS_WRITE, 2), 	-- 329
is_word(IS_READ, 764), 	-- 330
is_word(IS_WRITE, 2), 	-- 331
is_word(IS_READ, 763), 	-- 332
is_word(IS_WRITE, 762), 	-- 333
is_word(IS_READ, 761), 	-- 334
is_word(IS_WRITE, 2), 	-- 335
is_word(IS_READ, 760), 	-- 336
is_word(IS_WRITE, 2), 	-- 337
is_word(IS_READ, 759), 	-- 338
is_word(IS_WRITE, 2), 	-- 339
is_word(IS_READ, 758), 	-- 340
is_word(IS_WRITE, 757), 	-- 341
is_word(IS_READ, 756), 	-- 342
is_word(IS_WRITE, 755), 	-- 343
is_word(IS_READ, 196), 	-- 344
is_word(IS_GTE, 754), 	-- 345
is_word(IS_BRANCH, 753), 	-- 346
is_word(IS_READ, 752), 	-- 347
is_word(IS_WRITE, 751), 	-- 348
is_word(IS_READ, 197), 	-- 349
is_word(IS_GTE, 750), 	-- 350
is_word(IS_BRANCH, 749), 	-- 351
is_word(IS_READ, 196), 	-- 352
is_word(IS_EQ, 748), 	-- 353
is_word(IS_BRANCH, 747), 	-- 354
is_word(IS_READ, 196), 	-- 355
is_word(IS_EQ, 746), 	-- 356
is_word(IS_BRANCH, 745), 	-- 357
is_word(IS_READ, 197), 	-- 358
is_word(IS_EQ, 744), 	-- 359
is_word(IS_BRANCH, 743), 	-- 360
is_word(IS_READ, 197), 	-- 361
is_word(IS_EQ, 742), 	-- 362
is_word(IS_BRANCH, 741), 	-- 363
is_word(IS_READ, 196), 	-- 364
is_word(IS_OR, 197), 	-- 365
is_word(IS_AND, 740), 	-- 366
is_word(IS_EQ, 739), 	-- 367
is_word(IS_BRANCH, 738), 	-- 368
is_word(IS_READ, 737), 	-- 369
is_word(IS_WRITE, 736), 	-- 370
is_word(IS_READ, 196), 	-- 371
is_word(IS_MUL, 735), 	-- 372
is_word(IS_ADD, 197), 	-- 373
is_word(IS_ADD, 734), 	-- 374
is_word(IS_WRITE, 733), 	-- 375
is_word(IS_READ, 732), 	-- 376
is_word(IS_WRITE, 2), 	-- 377
is_word(IS_READ, 192), 	-- 378
is_word(IS_WRITE, 2), 	-- 379
is_word(IS_READ, 731), 	-- 380
is_word(IS_WRITE, 2), 	-- 381
is_word(IS_READ, 730), 	-- 382
is_word(IS_WRITE, 729), 	-- 383
is_word(IS_READ, 197), 	-- 384
is_word(IS_ADD, 728), 	-- 385
is_word(IS_WRITE, 727), 	-- 386
is_word(IS_READ, 726), 	-- 387
is_word(IS_WRITE, 725), 	-- 388
is_word(IS_READ, 196), 	-- 389
is_word(IS_ADD, 724), 	-- 390
is_word(IS_WRITE, 723), 	-- 391
is_word(IS_READ, 722), 	-- 392
is_word(IS_WRITE, 721), 	-- 393
is_word(IS_READ, 720), 	-- 394
is_word(IS_WRITE, 719), 	-- 395
is_word(IS_READ, 196), 	-- 396
is_word(IS_GTE, 718), 	-- 397
is_word(IS_BRANCH, 717), 	-- 398
is_word(IS_READ, 3), 	-- 399
is_word(IS_AND, 716), 	-- 400
is_word(IS_WRITE, 715), 	-- 401
is_word(IS_READ, 714), 	-- 402
is_word(IS_WRITE, 2), 	-- 403
is_word(IS_READ, 197), 	-- 404
is_word(IS_WRITE, 2), 	-- 405
is_word(IS_READ, 713), 	-- 406
is_word(IS_WRITE, 2), 	-- 407
is_word(IS_READ, 196), 	-- 408
is_word(IS_WRITE, 2), 	-- 409
is_word(IS_READ, 712), 	-- 410
is_word(IS_WRITE, 711), 	-- 411
is_word(IS_READ, 248), 	-- 412
is_word(IS_BRANCH, 710), 	-- 413
is_word(IS_READ, 196), 	-- 414
is_word(IS_ADD, 709), 	-- 415
is_word(IS_WRITE, 708), 	-- 416
is_word(IS_READ, 707), 	-- 417
is_word(IS_WRITE, 706), 	-- 418
is_word(IS_READ, 705), 	-- 419
is_word(IS_WRITE, 704), 	-- 420
is_word(IS_READ, 196), 	-- 421
is_word(IS_GTE, 703), 	-- 422
is_word(IS_BRANCH, 702), 	-- 423
is_word(IS_READ, 701), 	-- 424
is_word(IS_WRITE, 700), 	-- 425
is_word(IS_READ, 197), 	-- 426
is_word(IS_GTE, 699), 	-- 427
is_word(IS_BRANCH, 698), 	-- 428
is_word(IS_READ, 3), 	-- 429
is_word(IS_AND, 697), 	-- 430
is_word(IS_WRITE, 696), 	-- 431
is_word(IS_EQ, 695), 	-- 432
is_word(IS_BRANCH, 694), 	-- 433
is_word(IS_READ, 693), 	-- 434
is_word(IS_WRITE, 2), 	-- 435
is_word(IS_READ, 192), 	-- 436
is_word(IS_WRITE, 2), 	-- 437
is_word(IS_READ, 196), 	-- 438
is_word(IS_WRITE, 2), 	-- 439
is_word(IS_READ, 197), 	-- 440
is_word(IS_WRITE, 2), 	-- 441
is_word(IS_READ, 692), 	-- 442
is_word(IS_WRITE, 691), 	-- 443
is_word(IS_READ, 248), 	-- 444
is_word(IS_BRANCH, 690), 	-- 445
is_word(IS_READ, 197), 	-- 446
is_word(IS_ADD, 689), 	-- 447
is_word(IS_WRITE, 688), 	-- 448
is_word(IS_READ, 687), 	-- 449
is_word(IS_WRITE, 686), 	-- 450
is_word(IS_READ, 196), 	-- 451
is_word(IS_ADD, 685), 	-- 452
is_word(IS_WRITE, 684), 	-- 453
is_word(IS_READ, 683), 	-- 454
is_word(IS_WRITE, 682), 	-- 455
is_word(IS_READ, 681), 	-- 456
is_word(IS_WRITE, 680), 	-- 457
is_word(IS_READ, 2), 	-- 458
is_word(IS_WRITE, 679), 	-- 459
is_word(IS_ADD, 3), 	-- 460
is_word(IS_WRITE, 678), 	-- 461
is_word(IS_READ, 2), 	-- 462
is_word(IS_WRITE, 677), 	-- 463
is_word(IS_ADD, 3), 	-- 464
is_word(IS_WRITE, 676), 	-- 465
is_word(IS_READ, 2), 	-- 466
is_word(IS_WRITE, 675), 	-- 467
is_word(IS_ADD, 3), 	-- 468
is_word(IS_WRITE, 674), 	-- 469
is_word(IS_READ, 251), 	-- 470
is_word(IS_MUL, 673), 	-- 471
is_word(IS_ADD, 250), 	-- 472
is_word(IS_ADD, 672), 	-- 473
is_word(IS_WRITE, 671), 	-- 474
is_word(IS_READ, 252), 	-- 475
is_word(IS_NEQ, 670), 	-- 476
is_word(IS_BRANCH, 669), 	-- 477
is_word(IS_READ, 249), 	-- 478
is_word(IS_SUB, 668), 	-- 479
is_word(IS_WRITE, 667), 	-- 480
is_word(IS_READ, 666), 	-- 481
is_word(IS_WRITE, 665), 	-- 482
is_word(IS_READ, 252), 	-- 483
is_word(IS_NEQ, 664), 	-- 484
is_word(IS_BRANCH, 663), 	-- 485
is_word(IS_READ, 249), 	-- 486
is_word(IS_ADD, 662), 	-- 487
is_word(IS_WRITE, 661), 	-- 488
is_word(IS_READ, 660), 	-- 489
is_word(IS_WRITE, 659), 	-- 490
is_word(IS_READ, 252), 	-- 491
is_word(IS_NEQ, 658), 	-- 492
is_word(IS_BRANCH, 657), 	-- 493
is_word(IS_READ, 249), 	-- 494
is_word(IS_SUB, 656), 	-- 495
is_word(IS_WRITE, 655), 	-- 496
is_word(IS_READ, 654), 	-- 497
is_word(IS_WRITE, 653), 	-- 498
is_word(IS_READ, 252), 	-- 499
is_word(IS_NEQ, 652), 	-- 500
is_word(IS_BRANCH, 651), 	-- 501
is_word(IS_READ, 249), 	-- 502
is_word(IS_ADD, 650), 	-- 503
is_word(IS_WRITE, 649), 	-- 504
is_word(IS_READ, 648), 	-- 505
is_word(IS_WRITE, 647), 	-- 506
is_word(IS_READ, 249), 	-- 507
is_word(IS_WRITE, 646), 	-- 508
is_word(IS_ADD, 3), 	-- 509
is_word(IS_WRITE, 645), 	-- 510
is_word(IS_READ, 644), 	-- 511
is_word(IS_WRITE, 2), 	-- 512
is_word(IS_READ, 249), 	-- 513
is_word(IS_WRITE, 2), 	-- 514
is_word(IS_READ, 643), 	-- 515
is_word(IS_WRITE, 2), 	-- 516
is_word(IS_READ, 642), 	-- 517
is_word(IS_WRITE, 641), 	-- 518
is_word(IS_READ, 2), 	-- 519
is_word(IS_WRITE, 640), 	-- 520
is_word(IS_ADD, 3), 	-- 521
is_word(IS_WRITE, 639), 	-- 522
is_word(IS_READ, 2), 	-- 523
is_word(IS_WRITE, 638), 	-- 524
is_word(IS_ADD, 3), 	-- 525
is_word(IS_WRITE, 637), 	-- 526
is_word(IS_READ, 253), 	-- 527
is_word(IS_EQ, 636), 	-- 528
is_word(IS_BRANCH, 635), 	-- 529
is_word(IS_READ, 253), 	-- 530
is_word(IS_SUB, 634), 	-- 531
is_word(IS_WRITE, 633), 	-- 532
is_word(IS_READ, 632), 	-- 533
is_word(IS_WRITE, 631), 	-- 534
is_word(IS_READ, 2), 	-- 535
is_word(IS_WRITE, 630), 	-- 536
is_word(IS_ADD, 3), 	-- 537
is_word(IS_WRITE, 629), 	-- 538
is_word(IS_READ, 2), 	-- 539
is_word(IS_WRITE, 628), 	-- 540
is_word(IS_ADD, 3), 	-- 541
is_word(IS_WRITE, 627), 	-- 542
is_word(IS_READ, 2), 	-- 543
is_word(IS_WRITE, 626), 	-- 544
is_word(IS_ADD, 3), 	-- 545
is_word(IS_WRITE, 625), 	-- 546
is_word(IS_READ, 254), 	-- 547
is_word(IS_WRITE, 624), 	-- 548
is_word(IS_ADD, 3), 	-- 549
is_word(IS_EQ, 623), 	-- 550
is_word(IS_BRANCH, 622), 	-- 551
is_word(IS_READ, 254), 	-- 552
is_word(IS_WRITE, 621), 	-- 553
is_word(IS_ADD, 3), 	-- 554
is_word(IS_WRITE, 255), 	-- 555
is_word(IS_READ, 254), 	-- 556
is_word(IS_ADD, 620), 	-- 557
is_word(IS_WRITE, 619), 	-- 558
is_word(IS_READ, 255), 	-- 559
is_word(IS_ADD, 618), 	-- 560
is_word(IS_WRITE, 617), 	-- 561
is_word(IS_READ, 616), 	-- 562
is_word(IS_WRITE, 2), 	-- 563
is_word(IS_READ, 615), 	-- 564
is_word(IS_WRITE, 2), 	-- 565
is_word(IS_READ, 614), 	-- 566
is_word(IS_WRITE, 613), 	-- 567
is_word(IS_READ, 612), 	-- 568
is_word(IS_WRITE, 611), 	-- 569
is_word(IS_READ, 2), 	-- 570
is_word(IS_WRITE, 610), 	-- 571
is_word(IS_ADD, 3), 	-- 572
is_word(IS_WRITE, 609), 	-- 573
0, 	-- 574
0, 	-- 575
0, 	-- 576
0, 	-- 577
0, 	-- 578
0, 	-- 579
0, 	-- 580
0, 	-- 581
0, 	-- 582
0, 	-- 583
0, 	-- 584
0, 	-- 585
0, 	-- 586
0, 	-- 587
0, 	-- 588
0, 	-- 589
0, 	-- 590
0, 	-- 591
0, 	-- 592
0, 	-- 593
0, 	-- 594
0, 	-- 595
0, 	-- 596
0, 	-- 597
0, 	-- 598
0, 	-- 599
0, 	-- 600
0, 	-- 601
0, 	-- 602
0, 	-- 603
0, 	-- 604
0, 	-- 605
0, 	-- 606
0, 	-- 607
0, 	-- 608
0, 	-- 609
572, 	-- 610
0, 	-- 611
547, 	-- 612
0, 	-- 613
523, 	-- 614
4096, 	-- 615
568, 	-- 616
255, 	-- 617
1, 	-- 618
254, 	-- 619
1, 	-- 620
554, 	-- 621
570, 	-- 622
0, 	-- 623
549, 	-- 624
255, 	-- 625
545, 	-- 626
254, 	-- 627
541, 	-- 628
0, 	-- 629
537, 	-- 630
0, 	-- 631
527, 	-- 632
253, 	-- 633
1, 	-- 634
535, 	-- 635
0, 	-- 636
253, 	-- 637
525, 	-- 638
0, 	-- 639
521, 	-- 640
0, 	-- 641
539, 	-- 642
326, 	-- 643
519, 	-- 644
248, 	-- 645
509, 	-- 646
0, 	-- 647
507, 	-- 648
249, 	-- 649
1, 	-- 650
507, 	-- 651
3, 	-- 652
0, 	-- 653
507, 	-- 654
249, 	-- 655
1, 	-- 656
499, 	-- 657
2, 	-- 658
0, 	-- 659
507, 	-- 660
249, 	-- 661
40, 	-- 662
491, 	-- 663
1, 	-- 664
0, 	-- 665
507, 	-- 666
249, 	-- 667
40, 	-- 668
483, 	-- 669
0, 	-- 670
249, 	-- 671
1104, 	-- 672
40, 	-- 673
252, 	-- 674
468, 	-- 675
251, 	-- 676
464, 	-- 677
250, 	-- 678
460, 	-- 679
0, 	-- 680
456, 	-- 681
0, 	-- 682
421, 	-- 683
196, 	-- 684
2, 	-- 685
0, 	-- 686
426, 	-- 687
197, 	-- 688
2, 	-- 689
429, 	-- 690
0, 	-- 691
458, 	-- 692
444, 	-- 693
429, 	-- 694
0, 	-- 695
192, 	-- 696
3, 	-- 697
451, 	-- 698
37, 	-- 699
197, 	-- 700
2, 	-- 701
456, 	-- 702
21, 	-- 703
196, 	-- 704
4, 	-- 705
0, 	-- 706
396, 	-- 707
196, 	-- 708
2, 	-- 709
399, 	-- 710
0, 	-- 711
458, 	-- 712
2, 	-- 713
412, 	-- 714
197, 	-- 715
3, 	-- 716
419, 	-- 717
37, 	-- 718
196, 	-- 719
2, 	-- 720
0, 	-- 721
344, 	-- 722
196, 	-- 723
1, 	-- 724
0, 	-- 725
349, 	-- 726
197, 	-- 727
1, 	-- 728
0, 	-- 729
539, 	-- 730
326, 	-- 731
384, 	-- 732
192, 	-- 733
1104, 	-- 734
40, 	-- 735
0, 	-- 736
384, 	-- 737
371, 	-- 738
0, 	-- 739
1, 	-- 740
371, 	-- 741
38, 	-- 742
371, 	-- 743
0, 	-- 744
371, 	-- 745
22, 	-- 746
371, 	-- 747
0, 	-- 748
389, 	-- 749
39, 	-- 750
197, 	-- 751
0, 	-- 752
394, 	-- 753
23, 	-- 754
196, 	-- 755
0, 	-- 756
0, 	-- 757
539, 	-- 758
290, 	-- 759
1024, 	-- 760
342, 	-- 761
0, 	-- 762
523, 	-- 763
65536, 	-- 764
334, 	-- 765
0, 	-- 766
328	-- 767
