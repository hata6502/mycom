library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity osrom is
    port (addr	:in std_logic_vector (12 downto 0);
          data  :out std_logic_vector (7 downto 0)
         );
end osrom;

architecture arch_osrom of osrom is
begin
  process (addr)
  begin
    case addr(12 downto 0) is
      --addrbits 13
      --databits 8
      --varname data
      --little-endian
      --start_of_rom      -- rom2vhdl output.  Thu Jul 07 23:17:25 2016
      when "0000000000000" =>  data <= "00000010";  -- 0 = 2
      when "0000000000001" =>  data <= "11100000";  -- 1 = E0
      when "0000000000010" =>  data <= "01111000";  -- 2 = 78
      when "0000000000011" =>  data <= "11011000";  -- 3 = D8
      when "0000000000100" =>  data <= "10100010";  -- 4 = A2
      when "0000000000101" =>  data <= "11111111";  -- 5 = FF
      when "0000000000110" =>  data <= "10011010";  -- 6 = 9A
      when "0000000000111" =>  data <= "10101001";  -- 7 = A9
      when "0000000001000" =>  data <= "00000001";  -- 8 = 1
      when "0000000001001" =>  data <= "10000101";  -- 9 = 85
      when "0000000001010" =>  data <= "00010000";  -- A = 10
      when "0000000001011" =>  data <= "10101001";  -- B = A9
      when "0000000001100" =>  data <= "00000000";  -- C = 0
      when "0000000001101" =>  data <= "10000101";  -- D = 85
      when "0000000001110" =>  data <= "00010001";  -- E = 11
      when "0000000001111" =>  data <= "10100101";  -- F = A5
      when "0000000010000" =>  data <= "00010000";  -- 10 = 10
      when "0000000010001" =>  data <= "11001001";  -- 11 = C9
      when "0000000010010" =>  data <= "00000000";  -- 12 = 0
      when "0000000010011" =>  data <= "11110000";  -- 13 = F0
      when "0000000010100" =>  data <= "11111010";  -- 14 = FA
      when "0000000010101" =>  data <= "10101001";  -- 15 = A9
      when "0000000010110" =>  data <= "00000000";  -- 16 = 0
      when "0000000010111" =>  data <= "10000101";  -- 17 = 85
      when "0000000011000" =>  data <= "00010000";  -- 18 = 10
      when "0000000011001" =>  data <= "10100101";  -- 19 = A5
      when "0000000011010" =>  data <= "00010001";  -- 1A = 11
      when "0000000011011" =>  data <= "01001010";  -- 1B = 4A
      when "0000000011100" =>  data <= "01001010";  -- 1C = 4A
      when "0000000011101" =>  data <= "01001010";  -- 1D = 4A
      when "0000000011110" =>  data <= "01001010";  -- 1E = 4A
      when "0000000011111" =>  data <= "00011000";  -- 1F = 18
      when "0000000100000" =>  data <= "01101001";  -- 20 = 69
      when "0000000100001" =>  data <= "00110000";  -- 21 = 30
      when "0000000100010" =>  data <= "10001101";  -- 22 = 8D
      when "0000000100011" =>  data <= "00000000";  -- 23 = 0
      when "0000000100100" =>  data <= "00010001";  -- 24 = 11
      when "0000000100101" =>  data <= "10100101";  -- 25 = A5
      when "0000000100110" =>  data <= "00010001";  -- 26 = 11
      when "0000000100111" =>  data <= "00101001";  -- 27 = 29
      when "0000000101000" =>  data <= "00001111";  -- 28 = F
      when "0000000101001" =>  data <= "00011000";  -- 29 = 18
      when "0000000101010" =>  data <= "01101001";  -- 2A = 69
      when "0000000101011" =>  data <= "00110000";  -- 2B = 30
      when "0000000101100" =>  data <= "10001101";  -- 2C = 8D
      when "0000000101101" =>  data <= "00000001";  -- 2D = 1
      when "0000000101110" =>  data <= "00010001";  -- 2E = 11
      when "0000000101111" =>  data <= "10100101";  -- 2F = A5
      when "0000000110000" =>  data <= "00010001";  -- 30 = 11
      when "0000000110001" =>  data <= "10000101";  -- 31 = 85
      when "0000000110010" =>  data <= "00000000";  -- 32 = 0
      when "0000000110011" =>  data <= "11100110";  -- 33 = E6
      when "0000000110100" =>  data <= "00010001";  -- 34 = 11
      when "0000000110101" =>  data <= "01001100";  -- 35 = 4C
      when "0000000110110" =>  data <= "00001111";  -- 36 = F
      when "0000000110111" =>  data <= "11100000";  -- 37 = E0
      when "0000000111000" =>  data <= "01001000";  -- 38 = 48
      when "0000000111001" =>  data <= "10001010";  -- 39 = 8A
      when "0000000111010" =>  data <= "01001000";  -- 3A = 48
      when "0000000111011" =>  data <= "10011000";  -- 3B = 98
      when "0000000111100" =>  data <= "01001000";  -- 3C = 48
      when "0000000111101" =>  data <= "10101001";  -- 3D = A9
      when "0000000111110" =>  data <= "00000001";  -- 3E = 1
      when "0000000111111" =>  data <= "10000101";  -- 3F = 85
      when "0000001000000" =>  data <= "00010000";  -- 40 = 10
      when "0000001000001" =>  data <= "01101000";  -- 41 = 68
      when "0000001000010" =>  data <= "10101000";  -- 42 = A8
      when "0000001000011" =>  data <= "01101000";  -- 43 = 68
      when "0000001000100" =>  data <= "10101010";  -- 44 = AA
      when "0000001000101" =>  data <= "01101000";  -- 45 = 68
      when "0000001000110" =>  data <= "01000000";  -- 46 = 40
      when "0000001000111" =>  data <= "11111111";  -- 47 = FF
      when "0000001001000" =>  data <= "11111111";  -- 48 = FF
      when "0000001001001" =>  data <= "11111111";  -- 49 = FF
      when "0000001001010" =>  data <= "11111111";  -- 4A = FF
      when "0000001001011" =>  data <= "11111111";  -- 4B = FF
      when "0000001001100" =>  data <= "11111111";  -- 4C = FF
      when "0000001001101" =>  data <= "11111111";  -- 4D = FF
      when "0000001001110" =>  data <= "11111111";  -- 4E = FF
      when "0000001001111" =>  data <= "11111111";  -- 4F = FF
      when "0000001010000" =>  data <= "11111111";  -- 50 = FF
      when "0000001010001" =>  data <= "11111111";  -- 51 = FF
      when "0000001010010" =>  data <= "11111111";  -- 52 = FF
      when "0000001010011" =>  data <= "11111111";  -- 53 = FF
      when "0000001010100" =>  data <= "11111111";  -- 54 = FF
      when "0000001010101" =>  data <= "11111111";  -- 55 = FF
      when "0000001010110" =>  data <= "11111111";  -- 56 = FF
      when "0000001010111" =>  data <= "11111111";  -- 57 = FF
      when "0000001011000" =>  data <= "11111111";  -- 58 = FF
      when "0000001011001" =>  data <= "11111111";  -- 59 = FF
      when "0000001011010" =>  data <= "11111111";  -- 5A = FF
      when "0000001011011" =>  data <= "11111111";  -- 5B = FF
      when "0000001011100" =>  data <= "11111111";  -- 5C = FF
      when "0000001011101" =>  data <= "11111111";  -- 5D = FF
      when "0000001011110" =>  data <= "11111111";  -- 5E = FF
      when "0000001011111" =>  data <= "11111111";  -- 5F = FF
      when "0000001100000" =>  data <= "11111111";  -- 60 = FF
      when "0000001100001" =>  data <= "11111111";  -- 61 = FF
      when "0000001100010" =>  data <= "11111111";  -- 62 = FF
      when "0000001100011" =>  data <= "11111111";  -- 63 = FF
      when "0000001100100" =>  data <= "11111111";  -- 64 = FF
      when "0000001100101" =>  data <= "11111111";  -- 65 = FF
      when "0000001100110" =>  data <= "11111111";  -- 66 = FF
      when "0000001100111" =>  data <= "11111111";  -- 67 = FF
      when "0000001101000" =>  data <= "11111111";  -- 68 = FF
      when "0000001101001" =>  data <= "11111111";  -- 69 = FF
      when "0000001101010" =>  data <= "11111111";  -- 6A = FF
      when "0000001101011" =>  data <= "11111111";  -- 6B = FF
      when "0000001101100" =>  data <= "11111111";  -- 6C = FF
      when "0000001101101" =>  data <= "11111111";  -- 6D = FF
      when "0000001101110" =>  data <= "11111111";  -- 6E = FF
      when "0000001101111" =>  data <= "11111111";  -- 6F = FF
      when "0000001110000" =>  data <= "11111111";  -- 70 = FF
      when "0000001110001" =>  data <= "11111111";  -- 71 = FF
      when "0000001110010" =>  data <= "11111111";  -- 72 = FF
      when "0000001110011" =>  data <= "11111111";  -- 73 = FF
      when "0000001110100" =>  data <= "11111111";  -- 74 = FF
      when "0000001110101" =>  data <= "11111111";  -- 75 = FF
      when "0000001110110" =>  data <= "11111111";  -- 76 = FF
      when "0000001110111" =>  data <= "11111111";  -- 77 = FF
      when "0000001111000" =>  data <= "11111111";  -- 78 = FF
      when "0000001111001" =>  data <= "11111111";  -- 79 = FF
      when "0000001111010" =>  data <= "11111111";  -- 7A = FF
      when "0000001111011" =>  data <= "11111111";  -- 7B = FF
      when "0000001111100" =>  data <= "11111111";  -- 7C = FF
      when "0000001111101" =>  data <= "11111111";  -- 7D = FF
      when "0000001111110" =>  data <= "11111111";  -- 7E = FF
      when "0000001111111" =>  data <= "11111111";  -- 7F = FF
      when "0000010000000" =>  data <= "11111111";  -- 80 = FF
      when "0000010000001" =>  data <= "11111111";  -- 81 = FF
      when "0000010000010" =>  data <= "11111111";  -- 82 = FF
      when "0000010000011" =>  data <= "11111111";  -- 83 = FF
      when "0000010000100" =>  data <= "11111111";  -- 84 = FF
      when "0000010000101" =>  data <= "11111111";  -- 85 = FF
      when "0000010000110" =>  data <= "11111111";  -- 86 = FF
      when "0000010000111" =>  data <= "11111111";  -- 87 = FF
      when "0000010001000" =>  data <= "11111111";  -- 88 = FF
      when "0000010001001" =>  data <= "11111111";  -- 89 = FF
      when "0000010001010" =>  data <= "11111111";  -- 8A = FF
      when "0000010001011" =>  data <= "11111111";  -- 8B = FF
      when "0000010001100" =>  data <= "11111111";  -- 8C = FF
      when "0000010001101" =>  data <= "11111111";  -- 8D = FF
      when "0000010001110" =>  data <= "11111111";  -- 8E = FF
      when "0000010001111" =>  data <= "11111111";  -- 8F = FF
      when "0000010010000" =>  data <= "11111111";  -- 90 = FF
      when "0000010010001" =>  data <= "11111111";  -- 91 = FF
      when "0000010010010" =>  data <= "11111111";  -- 92 = FF
      when "0000010010011" =>  data <= "11111111";  -- 93 = FF
      when "0000010010100" =>  data <= "11111111";  -- 94 = FF
      when "0000010010101" =>  data <= "11111111";  -- 95 = FF
      when "0000010010110" =>  data <= "11111111";  -- 96 = FF
      when "0000010010111" =>  data <= "11111111";  -- 97 = FF
      when "0000010011000" =>  data <= "11111111";  -- 98 = FF
      when "0000010011001" =>  data <= "11111111";  -- 99 = FF
      when "0000010011010" =>  data <= "11111111";  -- 9A = FF
      when "0000010011011" =>  data <= "11111111";  -- 9B = FF
      when "0000010011100" =>  data <= "11111111";  -- 9C = FF
      when "0000010011101" =>  data <= "11111111";  -- 9D = FF
      when "0000010011110" =>  data <= "11111111";  -- 9E = FF
      when "0000010011111" =>  data <= "11111111";  -- 9F = FF
      when "0000010100000" =>  data <= "11111111";  -- A0 = FF
      when "0000010100001" =>  data <= "11111111";  -- A1 = FF
      when "0000010100010" =>  data <= "11111111";  -- A2 = FF
      when "0000010100011" =>  data <= "11111111";  -- A3 = FF
      when "0000010100100" =>  data <= "11111111";  -- A4 = FF
      when "0000010100101" =>  data <= "11111111";  -- A5 = FF
      when "0000010100110" =>  data <= "11111111";  -- A6 = FF
      when "0000010100111" =>  data <= "11111111";  -- A7 = FF
      when "0000010101000" =>  data <= "11111111";  -- A8 = FF
      when "0000010101001" =>  data <= "11111111";  -- A9 = FF
      when "0000010101010" =>  data <= "11111111";  -- AA = FF
      when "0000010101011" =>  data <= "11111111";  -- AB = FF
      when "0000010101100" =>  data <= "11111111";  -- AC = FF
      when "0000010101101" =>  data <= "11111111";  -- AD = FF
      when "0000010101110" =>  data <= "11111111";  -- AE = FF
      when "0000010101111" =>  data <= "11111111";  -- AF = FF
      when "0000010110000" =>  data <= "11111111";  -- B0 = FF
      when "0000010110001" =>  data <= "11111111";  -- B1 = FF
      when "0000010110010" =>  data <= "11111111";  -- B2 = FF
      when "0000010110011" =>  data <= "11111111";  -- B3 = FF
      when "0000010110100" =>  data <= "11111111";  -- B4 = FF
      when "0000010110101" =>  data <= "11111111";  -- B5 = FF
      when "0000010110110" =>  data <= "11111111";  -- B6 = FF
      when "0000010110111" =>  data <= "11111111";  -- B7 = FF
      when "0000010111000" =>  data <= "11111111";  -- B8 = FF
      when "0000010111001" =>  data <= "11111111";  -- B9 = FF
      when "0000010111010" =>  data <= "11111111";  -- BA = FF
      when "0000010111011" =>  data <= "11111111";  -- BB = FF
      when "0000010111100" =>  data <= "11111111";  -- BC = FF
      when "0000010111101" =>  data <= "11111111";  -- BD = FF
      when "0000010111110" =>  data <= "11111111";  -- BE = FF
      when "0000010111111" =>  data <= "11111111";  -- BF = FF
      when "0000011000000" =>  data <= "11111111";  -- C0 = FF
      when "0000011000001" =>  data <= "11111111";  -- C1 = FF
      when "0000011000010" =>  data <= "11111111";  -- C2 = FF
      when "0000011000011" =>  data <= "11111111";  -- C3 = FF
      when "0000011000100" =>  data <= "11111111";  -- C4 = FF
      when "0000011000101" =>  data <= "11111111";  -- C5 = FF
      when "0000011000110" =>  data <= "11111111";  -- C6 = FF
      when "0000011000111" =>  data <= "11111111";  -- C7 = FF
      when "0000011001000" =>  data <= "11111111";  -- C8 = FF
      when "0000011001001" =>  data <= "11111111";  -- C9 = FF
      when "0000011001010" =>  data <= "11111111";  -- CA = FF
      when "0000011001011" =>  data <= "11111111";  -- CB = FF
      when "0000011001100" =>  data <= "11111111";  -- CC = FF
      when "0000011001101" =>  data <= "11111111";  -- CD = FF
      when "0000011001110" =>  data <= "11111111";  -- CE = FF
      when "0000011001111" =>  data <= "11111111";  -- CF = FF
      when "0000011010000" =>  data <= "11111111";  -- D0 = FF
      when "0000011010001" =>  data <= "11111111";  -- D1 = FF
      when "0000011010010" =>  data <= "11111111";  -- D2 = FF
      when "0000011010011" =>  data <= "11111111";  -- D3 = FF
      when "0000011010100" =>  data <= "11111111";  -- D4 = FF
      when "0000011010101" =>  data <= "11111111";  -- D5 = FF
      when "0000011010110" =>  data <= "11111111";  -- D6 = FF
      when "0000011010111" =>  data <= "11111111";  -- D7 = FF
      when "0000011011000" =>  data <= "11111111";  -- D8 = FF
      when "0000011011001" =>  data <= "11111111";  -- D9 = FF
      when "0000011011010" =>  data <= "11111111";  -- DA = FF
      when "0000011011011" =>  data <= "11111111";  -- DB = FF
      when "0000011011100" =>  data <= "11111111";  -- DC = FF
      when "0000011011101" =>  data <= "11111111";  -- DD = FF
      when "0000011011110" =>  data <= "11111111";  -- DE = FF
      when "0000011011111" =>  data <= "11111111";  -- DF = FF
      when "0000011100000" =>  data <= "11111111";  -- E0 = FF
      when "0000011100001" =>  data <= "11111111";  -- E1 = FF
      when "0000011100010" =>  data <= "11111111";  -- E2 = FF
      when "0000011100011" =>  data <= "11111111";  -- E3 = FF
      when "0000011100100" =>  data <= "11111111";  -- E4 = FF
      when "0000011100101" =>  data <= "11111111";  -- E5 = FF
      when "0000011100110" =>  data <= "11111111";  -- E6 = FF
      when "0000011100111" =>  data <= "11111111";  -- E7 = FF
      when "0000011101000" =>  data <= "11111111";  -- E8 = FF
      when "0000011101001" =>  data <= "11111111";  -- E9 = FF
      when "0000011101010" =>  data <= "11111111";  -- EA = FF
      when "0000011101011" =>  data <= "11111111";  -- EB = FF
      when "0000011101100" =>  data <= "11111111";  -- EC = FF
      when "0000011101101" =>  data <= "11111111";  -- ED = FF
      when "0000011101110" =>  data <= "11111111";  -- EE = FF
      when "0000011101111" =>  data <= "11111111";  -- EF = FF
      when "0000011110000" =>  data <= "11111111";  -- F0 = FF
      when "0000011110001" =>  data <= "11111111";  -- F1 = FF
      when "0000011110010" =>  data <= "11111111";  -- F2 = FF
      when "0000011110011" =>  data <= "11111111";  -- F3 = FF
      when "0000011110100" =>  data <= "11111111";  -- F4 = FF
      when "0000011110101" =>  data <= "11111111";  -- F5 = FF
      when "0000011110110" =>  data <= "11111111";  -- F6 = FF
      when "0000011110111" =>  data <= "11111111";  -- F7 = FF
      when "0000011111000" =>  data <= "11111111";  -- F8 = FF
      when "0000011111001" =>  data <= "11111111";  -- F9 = FF
      when "0000011111010" =>  data <= "11111111";  -- FA = FF
      when "0000011111011" =>  data <= "11111111";  -- FB = FF
      when "0000011111100" =>  data <= "11111111";  -- FC = FF
      when "0000011111101" =>  data <= "11111111";  -- FD = FF
      when "0000011111110" =>  data <= "11111111";  -- FE = FF
      when "0000011111111" =>  data <= "11111111";  -- FF = FF
      when "0000100000000" =>  data <= "11111111";  -- 100 = FF
      when "0000100000001" =>  data <= "11111111";  -- 101 = FF
      when "0000100000010" =>  data <= "11111111";  -- 102 = FF
      when "0000100000011" =>  data <= "11111111";  -- 103 = FF
      when "0000100000100" =>  data <= "11111111";  -- 104 = FF
      when "0000100000101" =>  data <= "11111111";  -- 105 = FF
      when "0000100000110" =>  data <= "11111111";  -- 106 = FF
      when "0000100000111" =>  data <= "11111111";  -- 107 = FF
      when "0000100001000" =>  data <= "11111111";  -- 108 = FF
      when "0000100001001" =>  data <= "11111111";  -- 109 = FF
      when "0000100001010" =>  data <= "11111111";  -- 10A = FF
      when "0000100001011" =>  data <= "11111111";  -- 10B = FF
      when "0000100001100" =>  data <= "11111111";  -- 10C = FF
      when "0000100001101" =>  data <= "11111111";  -- 10D = FF
      when "0000100001110" =>  data <= "11111111";  -- 10E = FF
      when "0000100001111" =>  data <= "11111111";  -- 10F = FF
      when "0000100010000" =>  data <= "11111111";  -- 110 = FF
      when "0000100010001" =>  data <= "11111111";  -- 111 = FF
      when "0000100010010" =>  data <= "11111111";  -- 112 = FF
      when "0000100010011" =>  data <= "11111111";  -- 113 = FF
      when "0000100010100" =>  data <= "11111111";  -- 114 = FF
      when "0000100010101" =>  data <= "11111111";  -- 115 = FF
      when "0000100010110" =>  data <= "11111111";  -- 116 = FF
      when "0000100010111" =>  data <= "11111111";  -- 117 = FF
      when "0000100011000" =>  data <= "11111111";  -- 118 = FF
      when "0000100011001" =>  data <= "11111111";  -- 119 = FF
      when "0000100011010" =>  data <= "11111111";  -- 11A = FF
      when "0000100011011" =>  data <= "11111111";  -- 11B = FF
      when "0000100011100" =>  data <= "11111111";  -- 11C = FF
      when "0000100011101" =>  data <= "11111111";  -- 11D = FF
      when "0000100011110" =>  data <= "11111111";  -- 11E = FF
      when "0000100011111" =>  data <= "11111111";  -- 11F = FF
      when "0000100100000" =>  data <= "11111111";  -- 120 = FF
      when "0000100100001" =>  data <= "11111111";  -- 121 = FF
      when "0000100100010" =>  data <= "11111111";  -- 122 = FF
      when "0000100100011" =>  data <= "11111111";  -- 123 = FF
      when "0000100100100" =>  data <= "11111111";  -- 124 = FF
      when "0000100100101" =>  data <= "11111111";  -- 125 = FF
      when "0000100100110" =>  data <= "11111111";  -- 126 = FF
      when "0000100100111" =>  data <= "11111111";  -- 127 = FF
      when "0000100101000" =>  data <= "11111111";  -- 128 = FF
      when "0000100101001" =>  data <= "11111111";  -- 129 = FF
      when "0000100101010" =>  data <= "11111111";  -- 12A = FF
      when "0000100101011" =>  data <= "11111111";  -- 12B = FF
      when "0000100101100" =>  data <= "11111111";  -- 12C = FF
      when "0000100101101" =>  data <= "11111111";  -- 12D = FF
      when "0000100101110" =>  data <= "11111111";  -- 12E = FF
      when "0000100101111" =>  data <= "11111111";  -- 12F = FF
      when "0000100110000" =>  data <= "11111111";  -- 130 = FF
      when "0000100110001" =>  data <= "11111111";  -- 131 = FF
      when "0000100110010" =>  data <= "11111111";  -- 132 = FF
      when "0000100110011" =>  data <= "11111111";  -- 133 = FF
      when "0000100110100" =>  data <= "11111111";  -- 134 = FF
      when "0000100110101" =>  data <= "11111111";  -- 135 = FF
      when "0000100110110" =>  data <= "11111111";  -- 136 = FF
      when "0000100110111" =>  data <= "11111111";  -- 137 = FF
      when "0000100111000" =>  data <= "11111111";  -- 138 = FF
      when "0000100111001" =>  data <= "11111111";  -- 139 = FF
      when "0000100111010" =>  data <= "11111111";  -- 13A = FF
      when "0000100111011" =>  data <= "11111111";  -- 13B = FF
      when "0000100111100" =>  data <= "11111111";  -- 13C = FF
      when "0000100111101" =>  data <= "11111111";  -- 13D = FF
      when "0000100111110" =>  data <= "11111111";  -- 13E = FF
      when "0000100111111" =>  data <= "11111111";  -- 13F = FF
      when "0000101000000" =>  data <= "11111111";  -- 140 = FF
      when "0000101000001" =>  data <= "11111111";  -- 141 = FF
      when "0000101000010" =>  data <= "11111111";  -- 142 = FF
      when "0000101000011" =>  data <= "11111111";  -- 143 = FF
      when "0000101000100" =>  data <= "11111111";  -- 144 = FF
      when "0000101000101" =>  data <= "11111111";  -- 145 = FF
      when "0000101000110" =>  data <= "11111111";  -- 146 = FF
      when "0000101000111" =>  data <= "11111111";  -- 147 = FF
      when "0000101001000" =>  data <= "11111111";  -- 148 = FF
      when "0000101001001" =>  data <= "11111111";  -- 149 = FF
      when "0000101001010" =>  data <= "11111111";  -- 14A = FF
      when "0000101001011" =>  data <= "11111111";  -- 14B = FF
      when "0000101001100" =>  data <= "11111111";  -- 14C = FF
      when "0000101001101" =>  data <= "11111111";  -- 14D = FF
      when "0000101001110" =>  data <= "11111111";  -- 14E = FF
      when "0000101001111" =>  data <= "11111111";  -- 14F = FF
      when "0000101010000" =>  data <= "11111111";  -- 150 = FF
      when "0000101010001" =>  data <= "11111111";  -- 151 = FF
      when "0000101010010" =>  data <= "11111111";  -- 152 = FF
      when "0000101010011" =>  data <= "11111111";  -- 153 = FF
      when "0000101010100" =>  data <= "11111111";  -- 154 = FF
      when "0000101010101" =>  data <= "11111111";  -- 155 = FF
      when "0000101010110" =>  data <= "11111111";  -- 156 = FF
      when "0000101010111" =>  data <= "11111111";  -- 157 = FF
      when "0000101011000" =>  data <= "11111111";  -- 158 = FF
      when "0000101011001" =>  data <= "11111111";  -- 159 = FF
      when "0000101011010" =>  data <= "11111111";  -- 15A = FF
      when "0000101011011" =>  data <= "11111111";  -- 15B = FF
      when "0000101011100" =>  data <= "11111111";  -- 15C = FF
      when "0000101011101" =>  data <= "11111111";  -- 15D = FF
      when "0000101011110" =>  data <= "11111111";  -- 15E = FF
      when "0000101011111" =>  data <= "11111111";  -- 15F = FF
      when "0000101100000" =>  data <= "11111111";  -- 160 = FF
      when "0000101100001" =>  data <= "11111111";  -- 161 = FF
      when "0000101100010" =>  data <= "11111111";  -- 162 = FF
      when "0000101100011" =>  data <= "11111111";  -- 163 = FF
      when "0000101100100" =>  data <= "11111111";  -- 164 = FF
      when "0000101100101" =>  data <= "11111111";  -- 165 = FF
      when "0000101100110" =>  data <= "11111111";  -- 166 = FF
      when "0000101100111" =>  data <= "11111111";  -- 167 = FF
      when "0000101101000" =>  data <= "11111111";  -- 168 = FF
      when "0000101101001" =>  data <= "11111111";  -- 169 = FF
      when "0000101101010" =>  data <= "11111111";  -- 16A = FF
      when "0000101101011" =>  data <= "11111111";  -- 16B = FF
      when "0000101101100" =>  data <= "11111111";  -- 16C = FF
      when "0000101101101" =>  data <= "11111111";  -- 16D = FF
      when "0000101101110" =>  data <= "11111111";  -- 16E = FF
      when "0000101101111" =>  data <= "11111111";  -- 16F = FF
      when "0000101110000" =>  data <= "11111111";  -- 170 = FF
      when "0000101110001" =>  data <= "11111111";  -- 171 = FF
      when "0000101110010" =>  data <= "11111111";  -- 172 = FF
      when "0000101110011" =>  data <= "11111111";  -- 173 = FF
      when "0000101110100" =>  data <= "11111111";  -- 174 = FF
      when "0000101110101" =>  data <= "11111111";  -- 175 = FF
      when "0000101110110" =>  data <= "11111111";  -- 176 = FF
      when "0000101110111" =>  data <= "11111111";  -- 177 = FF
      when "0000101111000" =>  data <= "11111111";  -- 178 = FF
      when "0000101111001" =>  data <= "11111111";  -- 179 = FF
      when "0000101111010" =>  data <= "11111111";  -- 17A = FF
      when "0000101111011" =>  data <= "11111111";  -- 17B = FF
      when "0000101111100" =>  data <= "11111111";  -- 17C = FF
      when "0000101111101" =>  data <= "11111111";  -- 17D = FF
      when "0000101111110" =>  data <= "11111111";  -- 17E = FF
      when "0000101111111" =>  data <= "11111111";  -- 17F = FF
      when "0000110000000" =>  data <= "11111111";  -- 180 = FF
      when "0000110000001" =>  data <= "11111111";  -- 181 = FF
      when "0000110000010" =>  data <= "11111111";  -- 182 = FF
      when "0000110000011" =>  data <= "11111111";  -- 183 = FF
      when "0000110000100" =>  data <= "11111111";  -- 184 = FF
      when "0000110000101" =>  data <= "11111111";  -- 185 = FF
      when "0000110000110" =>  data <= "11111111";  -- 186 = FF
      when "0000110000111" =>  data <= "11111111";  -- 187 = FF
      when "0000110001000" =>  data <= "11111111";  -- 188 = FF
      when "0000110001001" =>  data <= "11111111";  -- 189 = FF
      when "0000110001010" =>  data <= "11111111";  -- 18A = FF
      when "0000110001011" =>  data <= "11111111";  -- 18B = FF
      when "0000110001100" =>  data <= "11111111";  -- 18C = FF
      when "0000110001101" =>  data <= "11111111";  -- 18D = FF
      when "0000110001110" =>  data <= "11111111";  -- 18E = FF
      when "0000110001111" =>  data <= "11111111";  -- 18F = FF
      when "0000110010000" =>  data <= "11111111";  -- 190 = FF
      when "0000110010001" =>  data <= "11111111";  -- 191 = FF
      when "0000110010010" =>  data <= "11111111";  -- 192 = FF
      when "0000110010011" =>  data <= "11111111";  -- 193 = FF
      when "0000110010100" =>  data <= "11111111";  -- 194 = FF
      when "0000110010101" =>  data <= "11111111";  -- 195 = FF
      when "0000110010110" =>  data <= "11111111";  -- 196 = FF
      when "0000110010111" =>  data <= "11111111";  -- 197 = FF
      when "0000110011000" =>  data <= "11111111";  -- 198 = FF
      when "0000110011001" =>  data <= "11111111";  -- 199 = FF
      when "0000110011010" =>  data <= "11111111";  -- 19A = FF
      when "0000110011011" =>  data <= "11111111";  -- 19B = FF
      when "0000110011100" =>  data <= "11111111";  -- 19C = FF
      when "0000110011101" =>  data <= "11111111";  -- 19D = FF
      when "0000110011110" =>  data <= "11111111";  -- 19E = FF
      when "0000110011111" =>  data <= "11111111";  -- 19F = FF
      when "0000110100000" =>  data <= "11111111";  -- 1A0 = FF
      when "0000110100001" =>  data <= "11111111";  -- 1A1 = FF
      when "0000110100010" =>  data <= "11111111";  -- 1A2 = FF
      when "0000110100011" =>  data <= "11111111";  -- 1A3 = FF
      when "0000110100100" =>  data <= "11111111";  -- 1A4 = FF
      when "0000110100101" =>  data <= "11111111";  -- 1A5 = FF
      when "0000110100110" =>  data <= "11111111";  -- 1A6 = FF
      when "0000110100111" =>  data <= "11111111";  -- 1A7 = FF
      when "0000110101000" =>  data <= "11111111";  -- 1A8 = FF
      when "0000110101001" =>  data <= "11111111";  -- 1A9 = FF
      when "0000110101010" =>  data <= "11111111";  -- 1AA = FF
      when "0000110101011" =>  data <= "11111111";  -- 1AB = FF
      when "0000110101100" =>  data <= "11111111";  -- 1AC = FF
      when "0000110101101" =>  data <= "11111111";  -- 1AD = FF
      when "0000110101110" =>  data <= "11111111";  -- 1AE = FF
      when "0000110101111" =>  data <= "11111111";  -- 1AF = FF
      when "0000110110000" =>  data <= "11111111";  -- 1B0 = FF
      when "0000110110001" =>  data <= "11111111";  -- 1B1 = FF
      when "0000110110010" =>  data <= "11111111";  -- 1B2 = FF
      when "0000110110011" =>  data <= "11111111";  -- 1B3 = FF
      when "0000110110100" =>  data <= "11111111";  -- 1B4 = FF
      when "0000110110101" =>  data <= "11111111";  -- 1B5 = FF
      when "0000110110110" =>  data <= "11111111";  -- 1B6 = FF
      when "0000110110111" =>  data <= "11111111";  -- 1B7 = FF
      when "0000110111000" =>  data <= "11111111";  -- 1B8 = FF
      when "0000110111001" =>  data <= "11111111";  -- 1B9 = FF
      when "0000110111010" =>  data <= "11111111";  -- 1BA = FF
      when "0000110111011" =>  data <= "11111111";  -- 1BB = FF
      when "0000110111100" =>  data <= "11111111";  -- 1BC = FF
      when "0000110111101" =>  data <= "11111111";  -- 1BD = FF
      when "0000110111110" =>  data <= "11111111";  -- 1BE = FF
      when "0000110111111" =>  data <= "11111111";  -- 1BF = FF
      when "0000111000000" =>  data <= "11111111";  -- 1C0 = FF
      when "0000111000001" =>  data <= "11111111";  -- 1C1 = FF
      when "0000111000010" =>  data <= "11111111";  -- 1C2 = FF
      when "0000111000011" =>  data <= "11111111";  -- 1C3 = FF
      when "0000111000100" =>  data <= "11111111";  -- 1C4 = FF
      when "0000111000101" =>  data <= "11111111";  -- 1C5 = FF
      when "0000111000110" =>  data <= "11111111";  -- 1C6 = FF
      when "0000111000111" =>  data <= "11111111";  -- 1C7 = FF
      when "0000111001000" =>  data <= "11111111";  -- 1C8 = FF
      when "0000111001001" =>  data <= "11111111";  -- 1C9 = FF
      when "0000111001010" =>  data <= "11111111";  -- 1CA = FF
      when "0000111001011" =>  data <= "11111111";  -- 1CB = FF
      when "0000111001100" =>  data <= "11111111";  -- 1CC = FF
      when "0000111001101" =>  data <= "11111111";  -- 1CD = FF
      when "0000111001110" =>  data <= "11111111";  -- 1CE = FF
      when "0000111001111" =>  data <= "11111111";  -- 1CF = FF
      when "0000111010000" =>  data <= "11111111";  -- 1D0 = FF
      when "0000111010001" =>  data <= "11111111";  -- 1D1 = FF
      when "0000111010010" =>  data <= "11111111";  -- 1D2 = FF
      when "0000111010011" =>  data <= "11111111";  -- 1D3 = FF
      when "0000111010100" =>  data <= "11111111";  -- 1D4 = FF
      when "0000111010101" =>  data <= "11111111";  -- 1D5 = FF
      when "0000111010110" =>  data <= "11111111";  -- 1D6 = FF
      when "0000111010111" =>  data <= "11111111";  -- 1D7 = FF
      when "0000111011000" =>  data <= "11111111";  -- 1D8 = FF
      when "0000111011001" =>  data <= "11111111";  -- 1D9 = FF
      when "0000111011010" =>  data <= "11111111";  -- 1DA = FF
      when "0000111011011" =>  data <= "11111111";  -- 1DB = FF
      when "0000111011100" =>  data <= "11111111";  -- 1DC = FF
      when "0000111011101" =>  data <= "11111111";  -- 1DD = FF
      when "0000111011110" =>  data <= "11111111";  -- 1DE = FF
      when "0000111011111" =>  data <= "11111111";  -- 1DF = FF
      when "0000111100000" =>  data <= "11111111";  -- 1E0 = FF
      when "0000111100001" =>  data <= "11111111";  -- 1E1 = FF
      when "0000111100010" =>  data <= "11111111";  -- 1E2 = FF
      when "0000111100011" =>  data <= "11111111";  -- 1E3 = FF
      when "0000111100100" =>  data <= "11111111";  -- 1E4 = FF
      when "0000111100101" =>  data <= "11111111";  -- 1E5 = FF
      when "0000111100110" =>  data <= "11111111";  -- 1E6 = FF
      when "0000111100111" =>  data <= "11111111";  -- 1E7 = FF
      when "0000111101000" =>  data <= "11111111";  -- 1E8 = FF
      when "0000111101001" =>  data <= "11111111";  -- 1E9 = FF
      when "0000111101010" =>  data <= "11111111";  -- 1EA = FF
      when "0000111101011" =>  data <= "11111111";  -- 1EB = FF
      when "0000111101100" =>  data <= "11111111";  -- 1EC = FF
      when "0000111101101" =>  data <= "11111111";  -- 1ED = FF
      when "0000111101110" =>  data <= "11111111";  -- 1EE = FF
      when "0000111101111" =>  data <= "11111111";  -- 1EF = FF
      when "0000111110000" =>  data <= "11111111";  -- 1F0 = FF
      when "0000111110001" =>  data <= "11111111";  -- 1F1 = FF
      when "0000111110010" =>  data <= "11111111";  -- 1F2 = FF
      when "0000111110011" =>  data <= "11111111";  -- 1F3 = FF
      when "0000111110100" =>  data <= "11111111";  -- 1F4 = FF
      when "0000111110101" =>  data <= "11111111";  -- 1F5 = FF
      when "0000111110110" =>  data <= "11111111";  -- 1F6 = FF
      when "0000111110111" =>  data <= "11111111";  -- 1F7 = FF
      when "0000111111000" =>  data <= "11111111";  -- 1F8 = FF
      when "0000111111001" =>  data <= "11111111";  -- 1F9 = FF
      when "0000111111010" =>  data <= "11111111";  -- 1FA = FF
      when "0000111111011" =>  data <= "11111111";  -- 1FB = FF
      when "0000111111100" =>  data <= "11111111";  -- 1FC = FF
      when "0000111111101" =>  data <= "11111111";  -- 1FD = FF
      when "0000111111110" =>  data <= "11111111";  -- 1FE = FF
      when "0000111111111" =>  data <= "11111111";  -- 1FF = FF
      when "0001000000000" =>  data <= "11111111";  -- 200 = FF
      when "0001000000001" =>  data <= "11111111";  -- 201 = FF
      when "0001000000010" =>  data <= "11111111";  -- 202 = FF
      when "0001000000011" =>  data <= "11111111";  -- 203 = FF
      when "0001000000100" =>  data <= "11111111";  -- 204 = FF
      when "0001000000101" =>  data <= "11111111";  -- 205 = FF
      when "0001000000110" =>  data <= "11111111";  -- 206 = FF
      when "0001000000111" =>  data <= "11111111";  -- 207 = FF
      when "0001000001000" =>  data <= "11111111";  -- 208 = FF
      when "0001000001001" =>  data <= "11111111";  -- 209 = FF
      when "0001000001010" =>  data <= "11111111";  -- 20A = FF
      when "0001000001011" =>  data <= "11111111";  -- 20B = FF
      when "0001000001100" =>  data <= "11111111";  -- 20C = FF
      when "0001000001101" =>  data <= "11111111";  -- 20D = FF
      when "0001000001110" =>  data <= "11111111";  -- 20E = FF
      when "0001000001111" =>  data <= "11111111";  -- 20F = FF
      when "0001000010000" =>  data <= "11111111";  -- 210 = FF
      when "0001000010001" =>  data <= "11111111";  -- 211 = FF
      when "0001000010010" =>  data <= "11111111";  -- 212 = FF
      when "0001000010011" =>  data <= "11111111";  -- 213 = FF
      when "0001000010100" =>  data <= "11111111";  -- 214 = FF
      when "0001000010101" =>  data <= "11111111";  -- 215 = FF
      when "0001000010110" =>  data <= "11111111";  -- 216 = FF
      when "0001000010111" =>  data <= "11111111";  -- 217 = FF
      when "0001000011000" =>  data <= "11111111";  -- 218 = FF
      when "0001000011001" =>  data <= "11111111";  -- 219 = FF
      when "0001000011010" =>  data <= "11111111";  -- 21A = FF
      when "0001000011011" =>  data <= "11111111";  -- 21B = FF
      when "0001000011100" =>  data <= "11111111";  -- 21C = FF
      when "0001000011101" =>  data <= "11111111";  -- 21D = FF
      when "0001000011110" =>  data <= "11111111";  -- 21E = FF
      when "0001000011111" =>  data <= "11111111";  -- 21F = FF
      when "0001000100000" =>  data <= "11111111";  -- 220 = FF
      when "0001000100001" =>  data <= "11111111";  -- 221 = FF
      when "0001000100010" =>  data <= "11111111";  -- 222 = FF
      when "0001000100011" =>  data <= "11111111";  -- 223 = FF
      when "0001000100100" =>  data <= "11111111";  -- 224 = FF
      when "0001000100101" =>  data <= "11111111";  -- 225 = FF
      when "0001000100110" =>  data <= "11111111";  -- 226 = FF
      when "0001000100111" =>  data <= "11111111";  -- 227 = FF
      when "0001000101000" =>  data <= "11111111";  -- 228 = FF
      when "0001000101001" =>  data <= "11111111";  -- 229 = FF
      when "0001000101010" =>  data <= "11111111";  -- 22A = FF
      when "0001000101011" =>  data <= "11111111";  -- 22B = FF
      when "0001000101100" =>  data <= "11111111";  -- 22C = FF
      when "0001000101101" =>  data <= "11111111";  -- 22D = FF
      when "0001000101110" =>  data <= "11111111";  -- 22E = FF
      when "0001000101111" =>  data <= "11111111";  -- 22F = FF
      when "0001000110000" =>  data <= "11111111";  -- 230 = FF
      when "0001000110001" =>  data <= "11111111";  -- 231 = FF
      when "0001000110010" =>  data <= "11111111";  -- 232 = FF
      when "0001000110011" =>  data <= "11111111";  -- 233 = FF
      when "0001000110100" =>  data <= "11111111";  -- 234 = FF
      when "0001000110101" =>  data <= "11111111";  -- 235 = FF
      when "0001000110110" =>  data <= "11111111";  -- 236 = FF
      when "0001000110111" =>  data <= "11111111";  -- 237 = FF
      when "0001000111000" =>  data <= "11111111";  -- 238 = FF
      when "0001000111001" =>  data <= "11111111";  -- 239 = FF
      when "0001000111010" =>  data <= "11111111";  -- 23A = FF
      when "0001000111011" =>  data <= "11111111";  -- 23B = FF
      when "0001000111100" =>  data <= "11111111";  -- 23C = FF
      when "0001000111101" =>  data <= "11111111";  -- 23D = FF
      when "0001000111110" =>  data <= "11111111";  -- 23E = FF
      when "0001000111111" =>  data <= "11111111";  -- 23F = FF
      when "0001001000000" =>  data <= "11111111";  -- 240 = FF
      when "0001001000001" =>  data <= "11111111";  -- 241 = FF
      when "0001001000010" =>  data <= "11111111";  -- 242 = FF
      when "0001001000011" =>  data <= "11111111";  -- 243 = FF
      when "0001001000100" =>  data <= "11111111";  -- 244 = FF
      when "0001001000101" =>  data <= "11111111";  -- 245 = FF
      when "0001001000110" =>  data <= "11111111";  -- 246 = FF
      when "0001001000111" =>  data <= "11111111";  -- 247 = FF
      when "0001001001000" =>  data <= "11111111";  -- 248 = FF
      when "0001001001001" =>  data <= "11111111";  -- 249 = FF
      when "0001001001010" =>  data <= "11111111";  -- 24A = FF
      when "0001001001011" =>  data <= "11111111";  -- 24B = FF
      when "0001001001100" =>  data <= "11111111";  -- 24C = FF
      when "0001001001101" =>  data <= "11111111";  -- 24D = FF
      when "0001001001110" =>  data <= "11111111";  -- 24E = FF
      when "0001001001111" =>  data <= "11111111";  -- 24F = FF
      when "0001001010000" =>  data <= "11111111";  -- 250 = FF
      when "0001001010001" =>  data <= "11111111";  -- 251 = FF
      when "0001001010010" =>  data <= "11111111";  -- 252 = FF
      when "0001001010011" =>  data <= "11111111";  -- 253 = FF
      when "0001001010100" =>  data <= "11111111";  -- 254 = FF
      when "0001001010101" =>  data <= "11111111";  -- 255 = FF
      when "0001001010110" =>  data <= "11111111";  -- 256 = FF
      when "0001001010111" =>  data <= "11111111";  -- 257 = FF
      when "0001001011000" =>  data <= "11111111";  -- 258 = FF
      when "0001001011001" =>  data <= "11111111";  -- 259 = FF
      when "0001001011010" =>  data <= "11111111";  -- 25A = FF
      when "0001001011011" =>  data <= "11111111";  -- 25B = FF
      when "0001001011100" =>  data <= "11111111";  -- 25C = FF
      when "0001001011101" =>  data <= "11111111";  -- 25D = FF
      when "0001001011110" =>  data <= "11111111";  -- 25E = FF
      when "0001001011111" =>  data <= "11111111";  -- 25F = FF
      when "0001001100000" =>  data <= "11111111";  -- 260 = FF
      when "0001001100001" =>  data <= "11111111";  -- 261 = FF
      when "0001001100010" =>  data <= "11111111";  -- 262 = FF
      when "0001001100011" =>  data <= "11111111";  -- 263 = FF
      when "0001001100100" =>  data <= "11111111";  -- 264 = FF
      when "0001001100101" =>  data <= "11111111";  -- 265 = FF
      when "0001001100110" =>  data <= "11111111";  -- 266 = FF
      when "0001001100111" =>  data <= "11111111";  -- 267 = FF
      when "0001001101000" =>  data <= "11111111";  -- 268 = FF
      when "0001001101001" =>  data <= "11111111";  -- 269 = FF
      when "0001001101010" =>  data <= "11111111";  -- 26A = FF
      when "0001001101011" =>  data <= "11111111";  -- 26B = FF
      when "0001001101100" =>  data <= "11111111";  -- 26C = FF
      when "0001001101101" =>  data <= "11111111";  -- 26D = FF
      when "0001001101110" =>  data <= "11111111";  -- 26E = FF
      when "0001001101111" =>  data <= "11111111";  -- 26F = FF
      when "0001001110000" =>  data <= "11111111";  -- 270 = FF
      when "0001001110001" =>  data <= "11111111";  -- 271 = FF
      when "0001001110010" =>  data <= "11111111";  -- 272 = FF
      when "0001001110011" =>  data <= "11111111";  -- 273 = FF
      when "0001001110100" =>  data <= "11111111";  -- 274 = FF
      when "0001001110101" =>  data <= "11111111";  -- 275 = FF
      when "0001001110110" =>  data <= "11111111";  -- 276 = FF
      when "0001001110111" =>  data <= "11111111";  -- 277 = FF
      when "0001001111000" =>  data <= "11111111";  -- 278 = FF
      when "0001001111001" =>  data <= "11111111";  -- 279 = FF
      when "0001001111010" =>  data <= "11111111";  -- 27A = FF
      when "0001001111011" =>  data <= "11111111";  -- 27B = FF
      when "0001001111100" =>  data <= "11111111";  -- 27C = FF
      when "0001001111101" =>  data <= "11111111";  -- 27D = FF
      when "0001001111110" =>  data <= "11111111";  -- 27E = FF
      when "0001001111111" =>  data <= "11111111";  -- 27F = FF
      when "0001010000000" =>  data <= "11111111";  -- 280 = FF
      when "0001010000001" =>  data <= "11111111";  -- 281 = FF
      when "0001010000010" =>  data <= "11111111";  -- 282 = FF
      when "0001010000011" =>  data <= "11111111";  -- 283 = FF
      when "0001010000100" =>  data <= "11111111";  -- 284 = FF
      when "0001010000101" =>  data <= "11111111";  -- 285 = FF
      when "0001010000110" =>  data <= "11111111";  -- 286 = FF
      when "0001010000111" =>  data <= "11111111";  -- 287 = FF
      when "0001010001000" =>  data <= "11111111";  -- 288 = FF
      when "0001010001001" =>  data <= "11111111";  -- 289 = FF
      when "0001010001010" =>  data <= "11111111";  -- 28A = FF
      when "0001010001011" =>  data <= "11111111";  -- 28B = FF
      when "0001010001100" =>  data <= "11111111";  -- 28C = FF
      when "0001010001101" =>  data <= "11111111";  -- 28D = FF
      when "0001010001110" =>  data <= "11111111";  -- 28E = FF
      when "0001010001111" =>  data <= "11111111";  -- 28F = FF
      when "0001010010000" =>  data <= "11111111";  -- 290 = FF
      when "0001010010001" =>  data <= "11111111";  -- 291 = FF
      when "0001010010010" =>  data <= "11111111";  -- 292 = FF
      when "0001010010011" =>  data <= "11111111";  -- 293 = FF
      when "0001010010100" =>  data <= "11111111";  -- 294 = FF
      when "0001010010101" =>  data <= "11111111";  -- 295 = FF
      when "0001010010110" =>  data <= "11111111";  -- 296 = FF
      when "0001010010111" =>  data <= "11111111";  -- 297 = FF
      when "0001010011000" =>  data <= "11111111";  -- 298 = FF
      when "0001010011001" =>  data <= "11111111";  -- 299 = FF
      when "0001010011010" =>  data <= "11111111";  -- 29A = FF
      when "0001010011011" =>  data <= "11111111";  -- 29B = FF
      when "0001010011100" =>  data <= "11111111";  -- 29C = FF
      when "0001010011101" =>  data <= "11111111";  -- 29D = FF
      when "0001010011110" =>  data <= "11111111";  -- 29E = FF
      when "0001010011111" =>  data <= "11111111";  -- 29F = FF
      when "0001010100000" =>  data <= "11111111";  -- 2A0 = FF
      when "0001010100001" =>  data <= "11111111";  -- 2A1 = FF
      when "0001010100010" =>  data <= "11111111";  -- 2A2 = FF
      when "0001010100011" =>  data <= "11111111";  -- 2A3 = FF
      when "0001010100100" =>  data <= "11111111";  -- 2A4 = FF
      when "0001010100101" =>  data <= "11111111";  -- 2A5 = FF
      when "0001010100110" =>  data <= "11111111";  -- 2A6 = FF
      when "0001010100111" =>  data <= "11111111";  -- 2A7 = FF
      when "0001010101000" =>  data <= "11111111";  -- 2A8 = FF
      when "0001010101001" =>  data <= "11111111";  -- 2A9 = FF
      when "0001010101010" =>  data <= "11111111";  -- 2AA = FF
      when "0001010101011" =>  data <= "11111111";  -- 2AB = FF
      when "0001010101100" =>  data <= "11111111";  -- 2AC = FF
      when "0001010101101" =>  data <= "11111111";  -- 2AD = FF
      when "0001010101110" =>  data <= "11111111";  -- 2AE = FF
      when "0001010101111" =>  data <= "11111111";  -- 2AF = FF
      when "0001010110000" =>  data <= "11111111";  -- 2B0 = FF
      when "0001010110001" =>  data <= "11111111";  -- 2B1 = FF
      when "0001010110010" =>  data <= "11111111";  -- 2B2 = FF
      when "0001010110011" =>  data <= "11111111";  -- 2B3 = FF
      when "0001010110100" =>  data <= "11111111";  -- 2B4 = FF
      when "0001010110101" =>  data <= "11111111";  -- 2B5 = FF
      when "0001010110110" =>  data <= "11111111";  -- 2B6 = FF
      when "0001010110111" =>  data <= "11111111";  -- 2B7 = FF
      when "0001010111000" =>  data <= "11111111";  -- 2B8 = FF
      when "0001010111001" =>  data <= "11111111";  -- 2B9 = FF
      when "0001010111010" =>  data <= "11111111";  -- 2BA = FF
      when "0001010111011" =>  data <= "11111111";  -- 2BB = FF
      when "0001010111100" =>  data <= "11111111";  -- 2BC = FF
      when "0001010111101" =>  data <= "11111111";  -- 2BD = FF
      when "0001010111110" =>  data <= "11111111";  -- 2BE = FF
      when "0001010111111" =>  data <= "11111111";  -- 2BF = FF
      when "0001011000000" =>  data <= "11111111";  -- 2C0 = FF
      when "0001011000001" =>  data <= "11111111";  -- 2C1 = FF
      when "0001011000010" =>  data <= "11111111";  -- 2C2 = FF
      when "0001011000011" =>  data <= "11111111";  -- 2C3 = FF
      when "0001011000100" =>  data <= "11111111";  -- 2C4 = FF
      when "0001011000101" =>  data <= "11111111";  -- 2C5 = FF
      when "0001011000110" =>  data <= "11111111";  -- 2C6 = FF
      when "0001011000111" =>  data <= "11111111";  -- 2C7 = FF
      when "0001011001000" =>  data <= "11111111";  -- 2C8 = FF
      when "0001011001001" =>  data <= "11111111";  -- 2C9 = FF
      when "0001011001010" =>  data <= "11111111";  -- 2CA = FF
      when "0001011001011" =>  data <= "11111111";  -- 2CB = FF
      when "0001011001100" =>  data <= "11111111";  -- 2CC = FF
      when "0001011001101" =>  data <= "11111111";  -- 2CD = FF
      when "0001011001110" =>  data <= "11111111";  -- 2CE = FF
      when "0001011001111" =>  data <= "11111111";  -- 2CF = FF
      when "0001011010000" =>  data <= "11111111";  -- 2D0 = FF
      when "0001011010001" =>  data <= "11111111";  -- 2D1 = FF
      when "0001011010010" =>  data <= "11111111";  -- 2D2 = FF
      when "0001011010011" =>  data <= "11111111";  -- 2D3 = FF
      when "0001011010100" =>  data <= "11111111";  -- 2D4 = FF
      when "0001011010101" =>  data <= "11111111";  -- 2D5 = FF
      when "0001011010110" =>  data <= "11111111";  -- 2D6 = FF
      when "0001011010111" =>  data <= "11111111";  -- 2D7 = FF
      when "0001011011000" =>  data <= "11111111";  -- 2D8 = FF
      when "0001011011001" =>  data <= "11111111";  -- 2D9 = FF
      when "0001011011010" =>  data <= "11111111";  -- 2DA = FF
      when "0001011011011" =>  data <= "11111111";  -- 2DB = FF
      when "0001011011100" =>  data <= "11111111";  -- 2DC = FF
      when "0001011011101" =>  data <= "11111111";  -- 2DD = FF
      when "0001011011110" =>  data <= "11111111";  -- 2DE = FF
      when "0001011011111" =>  data <= "11111111";  -- 2DF = FF
      when "0001011100000" =>  data <= "11111111";  -- 2E0 = FF
      when "0001011100001" =>  data <= "11111111";  -- 2E1 = FF
      when "0001011100010" =>  data <= "11111111";  -- 2E2 = FF
      when "0001011100011" =>  data <= "11111111";  -- 2E3 = FF
      when "0001011100100" =>  data <= "11111111";  -- 2E4 = FF
      when "0001011100101" =>  data <= "11111111";  -- 2E5 = FF
      when "0001011100110" =>  data <= "11111111";  -- 2E6 = FF
      when "0001011100111" =>  data <= "11111111";  -- 2E7 = FF
      when "0001011101000" =>  data <= "11111111";  -- 2E8 = FF
      when "0001011101001" =>  data <= "11111111";  -- 2E9 = FF
      when "0001011101010" =>  data <= "11111111";  -- 2EA = FF
      when "0001011101011" =>  data <= "11111111";  -- 2EB = FF
      when "0001011101100" =>  data <= "11111111";  -- 2EC = FF
      when "0001011101101" =>  data <= "11111111";  -- 2ED = FF
      when "0001011101110" =>  data <= "11111111";  -- 2EE = FF
      when "0001011101111" =>  data <= "11111111";  -- 2EF = FF
      when "0001011110000" =>  data <= "11111111";  -- 2F0 = FF
      when "0001011110001" =>  data <= "11111111";  -- 2F1 = FF
      when "0001011110010" =>  data <= "11111111";  -- 2F2 = FF
      when "0001011110011" =>  data <= "11111111";  -- 2F3 = FF
      when "0001011110100" =>  data <= "11111111";  -- 2F4 = FF
      when "0001011110101" =>  data <= "11111111";  -- 2F5 = FF
      when "0001011110110" =>  data <= "11111111";  -- 2F6 = FF
      when "0001011110111" =>  data <= "11111111";  -- 2F7 = FF
      when "0001011111000" =>  data <= "11111111";  -- 2F8 = FF
      when "0001011111001" =>  data <= "11111111";  -- 2F9 = FF
      when "0001011111010" =>  data <= "11111111";  -- 2FA = FF
      when "0001011111011" =>  data <= "11111111";  -- 2FB = FF
      when "0001011111100" =>  data <= "11111111";  -- 2FC = FF
      when "0001011111101" =>  data <= "11111111";  -- 2FD = FF
      when "0001011111110" =>  data <= "11111111";  -- 2FE = FF
      when "0001011111111" =>  data <= "11111111";  -- 2FF = FF
      when "0001100000000" =>  data <= "11111111";  -- 300 = FF
      when "0001100000001" =>  data <= "11111111";  -- 301 = FF
      when "0001100000010" =>  data <= "11111111";  -- 302 = FF
      when "0001100000011" =>  data <= "11111111";  -- 303 = FF
      when "0001100000100" =>  data <= "11111111";  -- 304 = FF
      when "0001100000101" =>  data <= "11111111";  -- 305 = FF
      when "0001100000110" =>  data <= "11111111";  -- 306 = FF
      when "0001100000111" =>  data <= "11111111";  -- 307 = FF
      when "0001100001000" =>  data <= "11111111";  -- 308 = FF
      when "0001100001001" =>  data <= "11111111";  -- 309 = FF
      when "0001100001010" =>  data <= "11111111";  -- 30A = FF
      when "0001100001011" =>  data <= "11111111";  -- 30B = FF
      when "0001100001100" =>  data <= "11111111";  -- 30C = FF
      when "0001100001101" =>  data <= "11111111";  -- 30D = FF
      when "0001100001110" =>  data <= "11111111";  -- 30E = FF
      when "0001100001111" =>  data <= "11111111";  -- 30F = FF
      when "0001100010000" =>  data <= "11111111";  -- 310 = FF
      when "0001100010001" =>  data <= "11111111";  -- 311 = FF
      when "0001100010010" =>  data <= "11111111";  -- 312 = FF
      when "0001100010011" =>  data <= "11111111";  -- 313 = FF
      when "0001100010100" =>  data <= "11111111";  -- 314 = FF
      when "0001100010101" =>  data <= "11111111";  -- 315 = FF
      when "0001100010110" =>  data <= "11111111";  -- 316 = FF
      when "0001100010111" =>  data <= "11111111";  -- 317 = FF
      when "0001100011000" =>  data <= "11111111";  -- 318 = FF
      when "0001100011001" =>  data <= "11111111";  -- 319 = FF
      when "0001100011010" =>  data <= "11111111";  -- 31A = FF
      when "0001100011011" =>  data <= "11111111";  -- 31B = FF
      when "0001100011100" =>  data <= "11111111";  -- 31C = FF
      when "0001100011101" =>  data <= "11111111";  -- 31D = FF
      when "0001100011110" =>  data <= "11111111";  -- 31E = FF
      when "0001100011111" =>  data <= "11111111";  -- 31F = FF
      when "0001100100000" =>  data <= "11111111";  -- 320 = FF
      when "0001100100001" =>  data <= "11111111";  -- 321 = FF
      when "0001100100010" =>  data <= "11111111";  -- 322 = FF
      when "0001100100011" =>  data <= "11111111";  -- 323 = FF
      when "0001100100100" =>  data <= "11111111";  -- 324 = FF
      when "0001100100101" =>  data <= "11111111";  -- 325 = FF
      when "0001100100110" =>  data <= "11111111";  -- 326 = FF
      when "0001100100111" =>  data <= "11111111";  -- 327 = FF
      when "0001100101000" =>  data <= "11111111";  -- 328 = FF
      when "0001100101001" =>  data <= "11111111";  -- 329 = FF
      when "0001100101010" =>  data <= "11111111";  -- 32A = FF
      when "0001100101011" =>  data <= "11111111";  -- 32B = FF
      when "0001100101100" =>  data <= "11111111";  -- 32C = FF
      when "0001100101101" =>  data <= "11111111";  -- 32D = FF
      when "0001100101110" =>  data <= "11111111";  -- 32E = FF
      when "0001100101111" =>  data <= "11111111";  -- 32F = FF
      when "0001100110000" =>  data <= "11111111";  -- 330 = FF
      when "0001100110001" =>  data <= "11111111";  -- 331 = FF
      when "0001100110010" =>  data <= "11111111";  -- 332 = FF
      when "0001100110011" =>  data <= "11111111";  -- 333 = FF
      when "0001100110100" =>  data <= "11111111";  -- 334 = FF
      when "0001100110101" =>  data <= "11111111";  -- 335 = FF
      when "0001100110110" =>  data <= "11111111";  -- 336 = FF
      when "0001100110111" =>  data <= "11111111";  -- 337 = FF
      when "0001100111000" =>  data <= "11111111";  -- 338 = FF
      when "0001100111001" =>  data <= "11111111";  -- 339 = FF
      when "0001100111010" =>  data <= "11111111";  -- 33A = FF
      when "0001100111011" =>  data <= "11111111";  -- 33B = FF
      when "0001100111100" =>  data <= "11111111";  -- 33C = FF
      when "0001100111101" =>  data <= "11111111";  -- 33D = FF
      when "0001100111110" =>  data <= "11111111";  -- 33E = FF
      when "0001100111111" =>  data <= "11111111";  -- 33F = FF
      when "0001101000000" =>  data <= "11111111";  -- 340 = FF
      when "0001101000001" =>  data <= "11111111";  -- 341 = FF
      when "0001101000010" =>  data <= "11111111";  -- 342 = FF
      when "0001101000011" =>  data <= "11111111";  -- 343 = FF
      when "0001101000100" =>  data <= "11111111";  -- 344 = FF
      when "0001101000101" =>  data <= "11111111";  -- 345 = FF
      when "0001101000110" =>  data <= "11111111";  -- 346 = FF
      when "0001101000111" =>  data <= "11111111";  -- 347 = FF
      when "0001101001000" =>  data <= "11111111";  -- 348 = FF
      when "0001101001001" =>  data <= "11111111";  -- 349 = FF
      when "0001101001010" =>  data <= "11111111";  -- 34A = FF
      when "0001101001011" =>  data <= "11111111";  -- 34B = FF
      when "0001101001100" =>  data <= "11111111";  -- 34C = FF
      when "0001101001101" =>  data <= "11111111";  -- 34D = FF
      when "0001101001110" =>  data <= "11111111";  -- 34E = FF
      when "0001101001111" =>  data <= "11111111";  -- 34F = FF
      when "0001101010000" =>  data <= "11111111";  -- 350 = FF
      when "0001101010001" =>  data <= "11111111";  -- 351 = FF
      when "0001101010010" =>  data <= "11111111";  -- 352 = FF
      when "0001101010011" =>  data <= "11111111";  -- 353 = FF
      when "0001101010100" =>  data <= "11111111";  -- 354 = FF
      when "0001101010101" =>  data <= "11111111";  -- 355 = FF
      when "0001101010110" =>  data <= "11111111";  -- 356 = FF
      when "0001101010111" =>  data <= "11111111";  -- 357 = FF
      when "0001101011000" =>  data <= "11111111";  -- 358 = FF
      when "0001101011001" =>  data <= "11111111";  -- 359 = FF
      when "0001101011010" =>  data <= "11111111";  -- 35A = FF
      when "0001101011011" =>  data <= "11111111";  -- 35B = FF
      when "0001101011100" =>  data <= "11111111";  -- 35C = FF
      when "0001101011101" =>  data <= "11111111";  -- 35D = FF
      when "0001101011110" =>  data <= "11111111";  -- 35E = FF
      when "0001101011111" =>  data <= "11111111";  -- 35F = FF
      when "0001101100000" =>  data <= "11111111";  -- 360 = FF
      when "0001101100001" =>  data <= "11111111";  -- 361 = FF
      when "0001101100010" =>  data <= "11111111";  -- 362 = FF
      when "0001101100011" =>  data <= "11111111";  -- 363 = FF
      when "0001101100100" =>  data <= "11111111";  -- 364 = FF
      when "0001101100101" =>  data <= "11111111";  -- 365 = FF
      when "0001101100110" =>  data <= "11111111";  -- 366 = FF
      when "0001101100111" =>  data <= "11111111";  -- 367 = FF
      when "0001101101000" =>  data <= "11111111";  -- 368 = FF
      when "0001101101001" =>  data <= "11111111";  -- 369 = FF
      when "0001101101010" =>  data <= "11111111";  -- 36A = FF
      when "0001101101011" =>  data <= "11111111";  -- 36B = FF
      when "0001101101100" =>  data <= "11111111";  -- 36C = FF
      when "0001101101101" =>  data <= "11111111";  -- 36D = FF
      when "0001101101110" =>  data <= "11111111";  -- 36E = FF
      when "0001101101111" =>  data <= "11111111";  -- 36F = FF
      when "0001101110000" =>  data <= "11111111";  -- 370 = FF
      when "0001101110001" =>  data <= "11111111";  -- 371 = FF
      when "0001101110010" =>  data <= "11111111";  -- 372 = FF
      when "0001101110011" =>  data <= "11111111";  -- 373 = FF
      when "0001101110100" =>  data <= "11111111";  -- 374 = FF
      when "0001101110101" =>  data <= "11111111";  -- 375 = FF
      when "0001101110110" =>  data <= "11111111";  -- 376 = FF
      when "0001101110111" =>  data <= "11111111";  -- 377 = FF
      when "0001101111000" =>  data <= "11111111";  -- 378 = FF
      when "0001101111001" =>  data <= "11111111";  -- 379 = FF
      when "0001101111010" =>  data <= "11111111";  -- 37A = FF
      when "0001101111011" =>  data <= "11111111";  -- 37B = FF
      when "0001101111100" =>  data <= "11111111";  -- 37C = FF
      when "0001101111101" =>  data <= "11111111";  -- 37D = FF
      when "0001101111110" =>  data <= "11111111";  -- 37E = FF
      when "0001101111111" =>  data <= "11111111";  -- 37F = FF
      when "0001110000000" =>  data <= "11111111";  -- 380 = FF
      when "0001110000001" =>  data <= "11111111";  -- 381 = FF
      when "0001110000010" =>  data <= "11111111";  -- 382 = FF
      when "0001110000011" =>  data <= "11111111";  -- 383 = FF
      when "0001110000100" =>  data <= "11111111";  -- 384 = FF
      when "0001110000101" =>  data <= "11111111";  -- 385 = FF
      when "0001110000110" =>  data <= "11111111";  -- 386 = FF
      when "0001110000111" =>  data <= "11111111";  -- 387 = FF
      when "0001110001000" =>  data <= "11111111";  -- 388 = FF
      when "0001110001001" =>  data <= "11111111";  -- 389 = FF
      when "0001110001010" =>  data <= "11111111";  -- 38A = FF
      when "0001110001011" =>  data <= "11111111";  -- 38B = FF
      when "0001110001100" =>  data <= "11111111";  -- 38C = FF
      when "0001110001101" =>  data <= "11111111";  -- 38D = FF
      when "0001110001110" =>  data <= "11111111";  -- 38E = FF
      when "0001110001111" =>  data <= "11111111";  -- 38F = FF
      when "0001110010000" =>  data <= "11111111";  -- 390 = FF
      when "0001110010001" =>  data <= "11111111";  -- 391 = FF
      when "0001110010010" =>  data <= "11111111";  -- 392 = FF
      when "0001110010011" =>  data <= "11111111";  -- 393 = FF
      when "0001110010100" =>  data <= "11111111";  -- 394 = FF
      when "0001110010101" =>  data <= "11111111";  -- 395 = FF
      when "0001110010110" =>  data <= "11111111";  -- 396 = FF
      when "0001110010111" =>  data <= "11111111";  -- 397 = FF
      when "0001110011000" =>  data <= "11111111";  -- 398 = FF
      when "0001110011001" =>  data <= "11111111";  -- 399 = FF
      when "0001110011010" =>  data <= "11111111";  -- 39A = FF
      when "0001110011011" =>  data <= "11111111";  -- 39B = FF
      when "0001110011100" =>  data <= "11111111";  -- 39C = FF
      when "0001110011101" =>  data <= "11111111";  -- 39D = FF
      when "0001110011110" =>  data <= "11111111";  -- 39E = FF
      when "0001110011111" =>  data <= "11111111";  -- 39F = FF
      when "0001110100000" =>  data <= "11111111";  -- 3A0 = FF
      when "0001110100001" =>  data <= "11111111";  -- 3A1 = FF
      when "0001110100010" =>  data <= "11111111";  -- 3A2 = FF
      when "0001110100011" =>  data <= "11111111";  -- 3A3 = FF
      when "0001110100100" =>  data <= "11111111";  -- 3A4 = FF
      when "0001110100101" =>  data <= "11111111";  -- 3A5 = FF
      when "0001110100110" =>  data <= "11111111";  -- 3A6 = FF
      when "0001110100111" =>  data <= "11111111";  -- 3A7 = FF
      when "0001110101000" =>  data <= "11111111";  -- 3A8 = FF
      when "0001110101001" =>  data <= "11111111";  -- 3A9 = FF
      when "0001110101010" =>  data <= "11111111";  -- 3AA = FF
      when "0001110101011" =>  data <= "11111111";  -- 3AB = FF
      when "0001110101100" =>  data <= "11111111";  -- 3AC = FF
      when "0001110101101" =>  data <= "11111111";  -- 3AD = FF
      when "0001110101110" =>  data <= "11111111";  -- 3AE = FF
      when "0001110101111" =>  data <= "11111111";  -- 3AF = FF
      when "0001110110000" =>  data <= "11111111";  -- 3B0 = FF
      when "0001110110001" =>  data <= "11111111";  -- 3B1 = FF
      when "0001110110010" =>  data <= "11111111";  -- 3B2 = FF
      when "0001110110011" =>  data <= "11111111";  -- 3B3 = FF
      when "0001110110100" =>  data <= "11111111";  -- 3B4 = FF
      when "0001110110101" =>  data <= "11111111";  -- 3B5 = FF
      when "0001110110110" =>  data <= "11111111";  -- 3B6 = FF
      when "0001110110111" =>  data <= "11111111";  -- 3B7 = FF
      when "0001110111000" =>  data <= "11111111";  -- 3B8 = FF
      when "0001110111001" =>  data <= "11111111";  -- 3B9 = FF
      when "0001110111010" =>  data <= "11111111";  -- 3BA = FF
      when "0001110111011" =>  data <= "11111111";  -- 3BB = FF
      when "0001110111100" =>  data <= "11111111";  -- 3BC = FF
      when "0001110111101" =>  data <= "11111111";  -- 3BD = FF
      when "0001110111110" =>  data <= "11111111";  -- 3BE = FF
      when "0001110111111" =>  data <= "11111111";  -- 3BF = FF
      when "0001111000000" =>  data <= "11111111";  -- 3C0 = FF
      when "0001111000001" =>  data <= "11111111";  -- 3C1 = FF
      when "0001111000010" =>  data <= "11111111";  -- 3C2 = FF
      when "0001111000011" =>  data <= "11111111";  -- 3C3 = FF
      when "0001111000100" =>  data <= "11111111";  -- 3C4 = FF
      when "0001111000101" =>  data <= "11111111";  -- 3C5 = FF
      when "0001111000110" =>  data <= "11111111";  -- 3C6 = FF
      when "0001111000111" =>  data <= "11111111";  -- 3C7 = FF
      when "0001111001000" =>  data <= "11111111";  -- 3C8 = FF
      when "0001111001001" =>  data <= "11111111";  -- 3C9 = FF
      when "0001111001010" =>  data <= "11111111";  -- 3CA = FF
      when "0001111001011" =>  data <= "11111111";  -- 3CB = FF
      when "0001111001100" =>  data <= "11111111";  -- 3CC = FF
      when "0001111001101" =>  data <= "11111111";  -- 3CD = FF
      when "0001111001110" =>  data <= "11111111";  -- 3CE = FF
      when "0001111001111" =>  data <= "11111111";  -- 3CF = FF
      when "0001111010000" =>  data <= "11111111";  -- 3D0 = FF
      when "0001111010001" =>  data <= "11111111";  -- 3D1 = FF
      when "0001111010010" =>  data <= "11111111";  -- 3D2 = FF
      when "0001111010011" =>  data <= "11111111";  -- 3D3 = FF
      when "0001111010100" =>  data <= "11111111";  -- 3D4 = FF
      when "0001111010101" =>  data <= "11111111";  -- 3D5 = FF
      when "0001111010110" =>  data <= "11111111";  -- 3D6 = FF
      when "0001111010111" =>  data <= "11111111";  -- 3D7 = FF
      when "0001111011000" =>  data <= "11111111";  -- 3D8 = FF
      when "0001111011001" =>  data <= "11111111";  -- 3D9 = FF
      when "0001111011010" =>  data <= "11111111";  -- 3DA = FF
      when "0001111011011" =>  data <= "11111111";  -- 3DB = FF
      when "0001111011100" =>  data <= "11111111";  -- 3DC = FF
      when "0001111011101" =>  data <= "11111111";  -- 3DD = FF
      when "0001111011110" =>  data <= "11111111";  -- 3DE = FF
      when "0001111011111" =>  data <= "11111111";  -- 3DF = FF
      when "0001111100000" =>  data <= "11111111";  -- 3E0 = FF
      when "0001111100001" =>  data <= "11111111";  -- 3E1 = FF
      when "0001111100010" =>  data <= "11111111";  -- 3E2 = FF
      when "0001111100011" =>  data <= "11111111";  -- 3E3 = FF
      when "0001111100100" =>  data <= "11111111";  -- 3E4 = FF
      when "0001111100101" =>  data <= "11111111";  -- 3E5 = FF
      when "0001111100110" =>  data <= "11111111";  -- 3E6 = FF
      when "0001111100111" =>  data <= "11111111";  -- 3E7 = FF
      when "0001111101000" =>  data <= "11111111";  -- 3E8 = FF
      when "0001111101001" =>  data <= "11111111";  -- 3E9 = FF
      when "0001111101010" =>  data <= "11111111";  -- 3EA = FF
      when "0001111101011" =>  data <= "11111111";  -- 3EB = FF
      when "0001111101100" =>  data <= "11111111";  -- 3EC = FF
      when "0001111101101" =>  data <= "11111111";  -- 3ED = FF
      when "0001111101110" =>  data <= "11111111";  -- 3EE = FF
      when "0001111101111" =>  data <= "11111111";  -- 3EF = FF
      when "0001111110000" =>  data <= "11111111";  -- 3F0 = FF
      when "0001111110001" =>  data <= "11111111";  -- 3F1 = FF
      when "0001111110010" =>  data <= "11111111";  -- 3F2 = FF
      when "0001111110011" =>  data <= "11111111";  -- 3F3 = FF
      when "0001111110100" =>  data <= "11111111";  -- 3F4 = FF
      when "0001111110101" =>  data <= "11111111";  -- 3F5 = FF
      when "0001111110110" =>  data <= "11111111";  -- 3F6 = FF
      when "0001111110111" =>  data <= "11111111";  -- 3F7 = FF
      when "0001111111000" =>  data <= "11111111";  -- 3F8 = FF
      when "0001111111001" =>  data <= "11111111";  -- 3F9 = FF
      when "0001111111010" =>  data <= "11111111";  -- 3FA = FF
      when "0001111111011" =>  data <= "11111111";  -- 3FB = FF
      when "0001111111100" =>  data <= "11111111";  -- 3FC = FF
      when "0001111111101" =>  data <= "11111111";  -- 3FD = FF
      when "0001111111110" =>  data <= "11111111";  -- 3FE = FF
      when "0001111111111" =>  data <= "11111111";  -- 3FF = FF
      when "0010000000000" =>  data <= "11111111";  -- 400 = FF
      when "0010000000001" =>  data <= "11111111";  -- 401 = FF
      when "0010000000010" =>  data <= "11111111";  -- 402 = FF
      when "0010000000011" =>  data <= "11111111";  -- 403 = FF
      when "0010000000100" =>  data <= "11111111";  -- 404 = FF
      when "0010000000101" =>  data <= "11111111";  -- 405 = FF
      when "0010000000110" =>  data <= "11111111";  -- 406 = FF
      when "0010000000111" =>  data <= "11111111";  -- 407 = FF
      when "0010000001000" =>  data <= "11111111";  -- 408 = FF
      when "0010000001001" =>  data <= "11111111";  -- 409 = FF
      when "0010000001010" =>  data <= "11111111";  -- 40A = FF
      when "0010000001011" =>  data <= "11111111";  -- 40B = FF
      when "0010000001100" =>  data <= "11111111";  -- 40C = FF
      when "0010000001101" =>  data <= "11111111";  -- 40D = FF
      when "0010000001110" =>  data <= "11111111";  -- 40E = FF
      when "0010000001111" =>  data <= "11111111";  -- 40F = FF
      when "0010000010000" =>  data <= "11111111";  -- 410 = FF
      when "0010000010001" =>  data <= "11111111";  -- 411 = FF
      when "0010000010010" =>  data <= "11111111";  -- 412 = FF
      when "0010000010011" =>  data <= "11111111";  -- 413 = FF
      when "0010000010100" =>  data <= "11111111";  -- 414 = FF
      when "0010000010101" =>  data <= "11111111";  -- 415 = FF
      when "0010000010110" =>  data <= "11111111";  -- 416 = FF
      when "0010000010111" =>  data <= "11111111";  -- 417 = FF
      when "0010000011000" =>  data <= "11111111";  -- 418 = FF
      when "0010000011001" =>  data <= "11111111";  -- 419 = FF
      when "0010000011010" =>  data <= "11111111";  -- 41A = FF
      when "0010000011011" =>  data <= "11111111";  -- 41B = FF
      when "0010000011100" =>  data <= "11111111";  -- 41C = FF
      when "0010000011101" =>  data <= "11111111";  -- 41D = FF
      when "0010000011110" =>  data <= "11111111";  -- 41E = FF
      when "0010000011111" =>  data <= "11111111";  -- 41F = FF
      when "0010000100000" =>  data <= "11111111";  -- 420 = FF
      when "0010000100001" =>  data <= "11111111";  -- 421 = FF
      when "0010000100010" =>  data <= "11111111";  -- 422 = FF
      when "0010000100011" =>  data <= "11111111";  -- 423 = FF
      when "0010000100100" =>  data <= "11111111";  -- 424 = FF
      when "0010000100101" =>  data <= "11111111";  -- 425 = FF
      when "0010000100110" =>  data <= "11111111";  -- 426 = FF
      when "0010000100111" =>  data <= "11111111";  -- 427 = FF
      when "0010000101000" =>  data <= "11111111";  -- 428 = FF
      when "0010000101001" =>  data <= "11111111";  -- 429 = FF
      when "0010000101010" =>  data <= "11111111";  -- 42A = FF
      when "0010000101011" =>  data <= "11111111";  -- 42B = FF
      when "0010000101100" =>  data <= "11111111";  -- 42C = FF
      when "0010000101101" =>  data <= "11111111";  -- 42D = FF
      when "0010000101110" =>  data <= "11111111";  -- 42E = FF
      when "0010000101111" =>  data <= "11111111";  -- 42F = FF
      when "0010000110000" =>  data <= "11111111";  -- 430 = FF
      when "0010000110001" =>  data <= "11111111";  -- 431 = FF
      when "0010000110010" =>  data <= "11111111";  -- 432 = FF
      when "0010000110011" =>  data <= "11111111";  -- 433 = FF
      when "0010000110100" =>  data <= "11111111";  -- 434 = FF
      when "0010000110101" =>  data <= "11111111";  -- 435 = FF
      when "0010000110110" =>  data <= "11111111";  -- 436 = FF
      when "0010000110111" =>  data <= "11111111";  -- 437 = FF
      when "0010000111000" =>  data <= "11111111";  -- 438 = FF
      when "0010000111001" =>  data <= "11111111";  -- 439 = FF
      when "0010000111010" =>  data <= "11111111";  -- 43A = FF
      when "0010000111011" =>  data <= "11111111";  -- 43B = FF
      when "0010000111100" =>  data <= "11111111";  -- 43C = FF
      when "0010000111101" =>  data <= "11111111";  -- 43D = FF
      when "0010000111110" =>  data <= "11111111";  -- 43E = FF
      when "0010000111111" =>  data <= "11111111";  -- 43F = FF
      when "0010001000000" =>  data <= "11111111";  -- 440 = FF
      when "0010001000001" =>  data <= "11111111";  -- 441 = FF
      when "0010001000010" =>  data <= "11111111";  -- 442 = FF
      when "0010001000011" =>  data <= "11111111";  -- 443 = FF
      when "0010001000100" =>  data <= "11111111";  -- 444 = FF
      when "0010001000101" =>  data <= "11111111";  -- 445 = FF
      when "0010001000110" =>  data <= "11111111";  -- 446 = FF
      when "0010001000111" =>  data <= "11111111";  -- 447 = FF
      when "0010001001000" =>  data <= "11111111";  -- 448 = FF
      when "0010001001001" =>  data <= "11111111";  -- 449 = FF
      when "0010001001010" =>  data <= "11111111";  -- 44A = FF
      when "0010001001011" =>  data <= "11111111";  -- 44B = FF
      when "0010001001100" =>  data <= "11111111";  -- 44C = FF
      when "0010001001101" =>  data <= "11111111";  -- 44D = FF
      when "0010001001110" =>  data <= "11111111";  -- 44E = FF
      when "0010001001111" =>  data <= "11111111";  -- 44F = FF
      when "0010001010000" =>  data <= "11111111";  -- 450 = FF
      when "0010001010001" =>  data <= "11111111";  -- 451 = FF
      when "0010001010010" =>  data <= "11111111";  -- 452 = FF
      when "0010001010011" =>  data <= "11111111";  -- 453 = FF
      when "0010001010100" =>  data <= "11111111";  -- 454 = FF
      when "0010001010101" =>  data <= "11111111";  -- 455 = FF
      when "0010001010110" =>  data <= "11111111";  -- 456 = FF
      when "0010001010111" =>  data <= "11111111";  -- 457 = FF
      when "0010001011000" =>  data <= "11111111";  -- 458 = FF
      when "0010001011001" =>  data <= "11111111";  -- 459 = FF
      when "0010001011010" =>  data <= "11111111";  -- 45A = FF
      when "0010001011011" =>  data <= "11111111";  -- 45B = FF
      when "0010001011100" =>  data <= "11111111";  -- 45C = FF
      when "0010001011101" =>  data <= "11111111";  -- 45D = FF
      when "0010001011110" =>  data <= "11111111";  -- 45E = FF
      when "0010001011111" =>  data <= "11111111";  -- 45F = FF
      when "0010001100000" =>  data <= "11111111";  -- 460 = FF
      when "0010001100001" =>  data <= "11111111";  -- 461 = FF
      when "0010001100010" =>  data <= "11111111";  -- 462 = FF
      when "0010001100011" =>  data <= "11111111";  -- 463 = FF
      when "0010001100100" =>  data <= "11111111";  -- 464 = FF
      when "0010001100101" =>  data <= "11111111";  -- 465 = FF
      when "0010001100110" =>  data <= "11111111";  -- 466 = FF
      when "0010001100111" =>  data <= "11111111";  -- 467 = FF
      when "0010001101000" =>  data <= "11111111";  -- 468 = FF
      when "0010001101001" =>  data <= "11111111";  -- 469 = FF
      when "0010001101010" =>  data <= "11111111";  -- 46A = FF
      when "0010001101011" =>  data <= "11111111";  -- 46B = FF
      when "0010001101100" =>  data <= "11111111";  -- 46C = FF
      when "0010001101101" =>  data <= "11111111";  -- 46D = FF
      when "0010001101110" =>  data <= "11111111";  -- 46E = FF
      when "0010001101111" =>  data <= "11111111";  -- 46F = FF
      when "0010001110000" =>  data <= "11111111";  -- 470 = FF
      when "0010001110001" =>  data <= "11111111";  -- 471 = FF
      when "0010001110010" =>  data <= "11111111";  -- 472 = FF
      when "0010001110011" =>  data <= "11111111";  -- 473 = FF
      when "0010001110100" =>  data <= "11111111";  -- 474 = FF
      when "0010001110101" =>  data <= "11111111";  -- 475 = FF
      when "0010001110110" =>  data <= "11111111";  -- 476 = FF
      when "0010001110111" =>  data <= "11111111";  -- 477 = FF
      when "0010001111000" =>  data <= "11111111";  -- 478 = FF
      when "0010001111001" =>  data <= "11111111";  -- 479 = FF
      when "0010001111010" =>  data <= "11111111";  -- 47A = FF
      when "0010001111011" =>  data <= "11111111";  -- 47B = FF
      when "0010001111100" =>  data <= "11111111";  -- 47C = FF
      when "0010001111101" =>  data <= "11111111";  -- 47D = FF
      when "0010001111110" =>  data <= "11111111";  -- 47E = FF
      when "0010001111111" =>  data <= "11111111";  -- 47F = FF
      when "0010010000000" =>  data <= "11111111";  -- 480 = FF
      when "0010010000001" =>  data <= "11111111";  -- 481 = FF
      when "0010010000010" =>  data <= "11111111";  -- 482 = FF
      when "0010010000011" =>  data <= "11111111";  -- 483 = FF
      when "0010010000100" =>  data <= "11111111";  -- 484 = FF
      when "0010010000101" =>  data <= "11111111";  -- 485 = FF
      when "0010010000110" =>  data <= "11111111";  -- 486 = FF
      when "0010010000111" =>  data <= "11111111";  -- 487 = FF
      when "0010010001000" =>  data <= "11111111";  -- 488 = FF
      when "0010010001001" =>  data <= "11111111";  -- 489 = FF
      when "0010010001010" =>  data <= "11111111";  -- 48A = FF
      when "0010010001011" =>  data <= "11111111";  -- 48B = FF
      when "0010010001100" =>  data <= "11111111";  -- 48C = FF
      when "0010010001101" =>  data <= "11111111";  -- 48D = FF
      when "0010010001110" =>  data <= "11111111";  -- 48E = FF
      when "0010010001111" =>  data <= "11111111";  -- 48F = FF
      when "0010010010000" =>  data <= "11111111";  -- 490 = FF
      when "0010010010001" =>  data <= "11111111";  -- 491 = FF
      when "0010010010010" =>  data <= "11111111";  -- 492 = FF
      when "0010010010011" =>  data <= "11111111";  -- 493 = FF
      when "0010010010100" =>  data <= "11111111";  -- 494 = FF
      when "0010010010101" =>  data <= "11111111";  -- 495 = FF
      when "0010010010110" =>  data <= "11111111";  -- 496 = FF
      when "0010010010111" =>  data <= "11111111";  -- 497 = FF
      when "0010010011000" =>  data <= "11111111";  -- 498 = FF
      when "0010010011001" =>  data <= "11111111";  -- 499 = FF
      when "0010010011010" =>  data <= "11111111";  -- 49A = FF
      when "0010010011011" =>  data <= "11111111";  -- 49B = FF
      when "0010010011100" =>  data <= "11111111";  -- 49C = FF
      when "0010010011101" =>  data <= "11111111";  -- 49D = FF
      when "0010010011110" =>  data <= "11111111";  -- 49E = FF
      when "0010010011111" =>  data <= "11111111";  -- 49F = FF
      when "0010010100000" =>  data <= "11111111";  -- 4A0 = FF
      when "0010010100001" =>  data <= "11111111";  -- 4A1 = FF
      when "0010010100010" =>  data <= "11111111";  -- 4A2 = FF
      when "0010010100011" =>  data <= "11111111";  -- 4A3 = FF
      when "0010010100100" =>  data <= "11111111";  -- 4A4 = FF
      when "0010010100101" =>  data <= "11111111";  -- 4A5 = FF
      when "0010010100110" =>  data <= "11111111";  -- 4A6 = FF
      when "0010010100111" =>  data <= "11111111";  -- 4A7 = FF
      when "0010010101000" =>  data <= "11111111";  -- 4A8 = FF
      when "0010010101001" =>  data <= "11111111";  -- 4A9 = FF
      when "0010010101010" =>  data <= "11111111";  -- 4AA = FF
      when "0010010101011" =>  data <= "11111111";  -- 4AB = FF
      when "0010010101100" =>  data <= "11111111";  -- 4AC = FF
      when "0010010101101" =>  data <= "11111111";  -- 4AD = FF
      when "0010010101110" =>  data <= "11111111";  -- 4AE = FF
      when "0010010101111" =>  data <= "11111111";  -- 4AF = FF
      when "0010010110000" =>  data <= "11111111";  -- 4B0 = FF
      when "0010010110001" =>  data <= "11111111";  -- 4B1 = FF
      when "0010010110010" =>  data <= "11111111";  -- 4B2 = FF
      when "0010010110011" =>  data <= "11111111";  -- 4B3 = FF
      when "0010010110100" =>  data <= "11111111";  -- 4B4 = FF
      when "0010010110101" =>  data <= "11111111";  -- 4B5 = FF
      when "0010010110110" =>  data <= "11111111";  -- 4B6 = FF
      when "0010010110111" =>  data <= "11111111";  -- 4B7 = FF
      when "0010010111000" =>  data <= "11111111";  -- 4B8 = FF
      when "0010010111001" =>  data <= "11111111";  -- 4B9 = FF
      when "0010010111010" =>  data <= "11111111";  -- 4BA = FF
      when "0010010111011" =>  data <= "11111111";  -- 4BB = FF
      when "0010010111100" =>  data <= "11111111";  -- 4BC = FF
      when "0010010111101" =>  data <= "11111111";  -- 4BD = FF
      when "0010010111110" =>  data <= "11111111";  -- 4BE = FF
      when "0010010111111" =>  data <= "11111111";  -- 4BF = FF
      when "0010011000000" =>  data <= "11111111";  -- 4C0 = FF
      when "0010011000001" =>  data <= "11111111";  -- 4C1 = FF
      when "0010011000010" =>  data <= "11111111";  -- 4C2 = FF
      when "0010011000011" =>  data <= "11111111";  -- 4C3 = FF
      when "0010011000100" =>  data <= "11111111";  -- 4C4 = FF
      when "0010011000101" =>  data <= "11111111";  -- 4C5 = FF
      when "0010011000110" =>  data <= "11111111";  -- 4C6 = FF
      when "0010011000111" =>  data <= "11111111";  -- 4C7 = FF
      when "0010011001000" =>  data <= "11111111";  -- 4C8 = FF
      when "0010011001001" =>  data <= "11111111";  -- 4C9 = FF
      when "0010011001010" =>  data <= "11111111";  -- 4CA = FF
      when "0010011001011" =>  data <= "11111111";  -- 4CB = FF
      when "0010011001100" =>  data <= "11111111";  -- 4CC = FF
      when "0010011001101" =>  data <= "11111111";  -- 4CD = FF
      when "0010011001110" =>  data <= "11111111";  -- 4CE = FF
      when "0010011001111" =>  data <= "11111111";  -- 4CF = FF
      when "0010011010000" =>  data <= "11111111";  -- 4D0 = FF
      when "0010011010001" =>  data <= "11111111";  -- 4D1 = FF
      when "0010011010010" =>  data <= "11111111";  -- 4D2 = FF
      when "0010011010011" =>  data <= "11111111";  -- 4D3 = FF
      when "0010011010100" =>  data <= "11111111";  -- 4D4 = FF
      when "0010011010101" =>  data <= "11111111";  -- 4D5 = FF
      when "0010011010110" =>  data <= "11111111";  -- 4D6 = FF
      when "0010011010111" =>  data <= "11111111";  -- 4D7 = FF
      when "0010011011000" =>  data <= "11111111";  -- 4D8 = FF
      when "0010011011001" =>  data <= "11111111";  -- 4D9 = FF
      when "0010011011010" =>  data <= "11111111";  -- 4DA = FF
      when "0010011011011" =>  data <= "11111111";  -- 4DB = FF
      when "0010011011100" =>  data <= "11111111";  -- 4DC = FF
      when "0010011011101" =>  data <= "11111111";  -- 4DD = FF
      when "0010011011110" =>  data <= "11111111";  -- 4DE = FF
      when "0010011011111" =>  data <= "11111111";  -- 4DF = FF
      when "0010011100000" =>  data <= "11111111";  -- 4E0 = FF
      when "0010011100001" =>  data <= "11111111";  -- 4E1 = FF
      when "0010011100010" =>  data <= "11111111";  -- 4E2 = FF
      when "0010011100011" =>  data <= "11111111";  -- 4E3 = FF
      when "0010011100100" =>  data <= "11111111";  -- 4E4 = FF
      when "0010011100101" =>  data <= "11111111";  -- 4E5 = FF
      when "0010011100110" =>  data <= "11111111";  -- 4E6 = FF
      when "0010011100111" =>  data <= "11111111";  -- 4E7 = FF
      when "0010011101000" =>  data <= "11111111";  -- 4E8 = FF
      when "0010011101001" =>  data <= "11111111";  -- 4E9 = FF
      when "0010011101010" =>  data <= "11111111";  -- 4EA = FF
      when "0010011101011" =>  data <= "11111111";  -- 4EB = FF
      when "0010011101100" =>  data <= "11111111";  -- 4EC = FF
      when "0010011101101" =>  data <= "11111111";  -- 4ED = FF
      when "0010011101110" =>  data <= "11111111";  -- 4EE = FF
      when "0010011101111" =>  data <= "11111111";  -- 4EF = FF
      when "0010011110000" =>  data <= "11111111";  -- 4F0 = FF
      when "0010011110001" =>  data <= "11111111";  -- 4F1 = FF
      when "0010011110010" =>  data <= "11111111";  -- 4F2 = FF
      when "0010011110011" =>  data <= "11111111";  -- 4F3 = FF
      when "0010011110100" =>  data <= "11111111";  -- 4F4 = FF
      when "0010011110101" =>  data <= "11111111";  -- 4F5 = FF
      when "0010011110110" =>  data <= "11111111";  -- 4F6 = FF
      when "0010011110111" =>  data <= "11111111";  -- 4F7 = FF
      when "0010011111000" =>  data <= "11111111";  -- 4F8 = FF
      when "0010011111001" =>  data <= "11111111";  -- 4F9 = FF
      when "0010011111010" =>  data <= "11111111";  -- 4FA = FF
      when "0010011111011" =>  data <= "11111111";  -- 4FB = FF
      when "0010011111100" =>  data <= "11111111";  -- 4FC = FF
      when "0010011111101" =>  data <= "11111111";  -- 4FD = FF
      when "0010011111110" =>  data <= "11111111";  -- 4FE = FF
      when "0010011111111" =>  data <= "11111111";  -- 4FF = FF
      when "0010100000000" =>  data <= "11111111";  -- 500 = FF
      when "0010100000001" =>  data <= "11111111";  -- 501 = FF
      when "0010100000010" =>  data <= "11111111";  -- 502 = FF
      when "0010100000011" =>  data <= "11111111";  -- 503 = FF
      when "0010100000100" =>  data <= "11111111";  -- 504 = FF
      when "0010100000101" =>  data <= "11111111";  -- 505 = FF
      when "0010100000110" =>  data <= "11111111";  -- 506 = FF
      when "0010100000111" =>  data <= "11111111";  -- 507 = FF
      when "0010100001000" =>  data <= "11111111";  -- 508 = FF
      when "0010100001001" =>  data <= "11111111";  -- 509 = FF
      when "0010100001010" =>  data <= "11111111";  -- 50A = FF
      when "0010100001011" =>  data <= "11111111";  -- 50B = FF
      when "0010100001100" =>  data <= "11111111";  -- 50C = FF
      when "0010100001101" =>  data <= "11111111";  -- 50D = FF
      when "0010100001110" =>  data <= "11111111";  -- 50E = FF
      when "0010100001111" =>  data <= "11111111";  -- 50F = FF
      when "0010100010000" =>  data <= "11111111";  -- 510 = FF
      when "0010100010001" =>  data <= "11111111";  -- 511 = FF
      when "0010100010010" =>  data <= "11111111";  -- 512 = FF
      when "0010100010011" =>  data <= "11111111";  -- 513 = FF
      when "0010100010100" =>  data <= "11111111";  -- 514 = FF
      when "0010100010101" =>  data <= "11111111";  -- 515 = FF
      when "0010100010110" =>  data <= "11111111";  -- 516 = FF
      when "0010100010111" =>  data <= "11111111";  -- 517 = FF
      when "0010100011000" =>  data <= "11111111";  -- 518 = FF
      when "0010100011001" =>  data <= "11111111";  -- 519 = FF
      when "0010100011010" =>  data <= "11111111";  -- 51A = FF
      when "0010100011011" =>  data <= "11111111";  -- 51B = FF
      when "0010100011100" =>  data <= "11111111";  -- 51C = FF
      when "0010100011101" =>  data <= "11111111";  -- 51D = FF
      when "0010100011110" =>  data <= "11111111";  -- 51E = FF
      when "0010100011111" =>  data <= "11111111";  -- 51F = FF
      when "0010100100000" =>  data <= "11111111";  -- 520 = FF
      when "0010100100001" =>  data <= "11111111";  -- 521 = FF
      when "0010100100010" =>  data <= "11111111";  -- 522 = FF
      when "0010100100011" =>  data <= "11111111";  -- 523 = FF
      when "0010100100100" =>  data <= "11111111";  -- 524 = FF
      when "0010100100101" =>  data <= "11111111";  -- 525 = FF
      when "0010100100110" =>  data <= "11111111";  -- 526 = FF
      when "0010100100111" =>  data <= "11111111";  -- 527 = FF
      when "0010100101000" =>  data <= "11111111";  -- 528 = FF
      when "0010100101001" =>  data <= "11111111";  -- 529 = FF
      when "0010100101010" =>  data <= "11111111";  -- 52A = FF
      when "0010100101011" =>  data <= "11111111";  -- 52B = FF
      when "0010100101100" =>  data <= "11111111";  -- 52C = FF
      when "0010100101101" =>  data <= "11111111";  -- 52D = FF
      when "0010100101110" =>  data <= "11111111";  -- 52E = FF
      when "0010100101111" =>  data <= "11111111";  -- 52F = FF
      when "0010100110000" =>  data <= "11111111";  -- 530 = FF
      when "0010100110001" =>  data <= "11111111";  -- 531 = FF
      when "0010100110010" =>  data <= "11111111";  -- 532 = FF
      when "0010100110011" =>  data <= "11111111";  -- 533 = FF
      when "0010100110100" =>  data <= "11111111";  -- 534 = FF
      when "0010100110101" =>  data <= "11111111";  -- 535 = FF
      when "0010100110110" =>  data <= "11111111";  -- 536 = FF
      when "0010100110111" =>  data <= "11111111";  -- 537 = FF
      when "0010100111000" =>  data <= "11111111";  -- 538 = FF
      when "0010100111001" =>  data <= "11111111";  -- 539 = FF
      when "0010100111010" =>  data <= "11111111";  -- 53A = FF
      when "0010100111011" =>  data <= "11111111";  -- 53B = FF
      when "0010100111100" =>  data <= "11111111";  -- 53C = FF
      when "0010100111101" =>  data <= "11111111";  -- 53D = FF
      when "0010100111110" =>  data <= "11111111";  -- 53E = FF
      when "0010100111111" =>  data <= "11111111";  -- 53F = FF
      when "0010101000000" =>  data <= "11111111";  -- 540 = FF
      when "0010101000001" =>  data <= "11111111";  -- 541 = FF
      when "0010101000010" =>  data <= "11111111";  -- 542 = FF
      when "0010101000011" =>  data <= "11111111";  -- 543 = FF
      when "0010101000100" =>  data <= "11111111";  -- 544 = FF
      when "0010101000101" =>  data <= "11111111";  -- 545 = FF
      when "0010101000110" =>  data <= "11111111";  -- 546 = FF
      when "0010101000111" =>  data <= "11111111";  -- 547 = FF
      when "0010101001000" =>  data <= "11111111";  -- 548 = FF
      when "0010101001001" =>  data <= "11111111";  -- 549 = FF
      when "0010101001010" =>  data <= "11111111";  -- 54A = FF
      when "0010101001011" =>  data <= "11111111";  -- 54B = FF
      when "0010101001100" =>  data <= "11111111";  -- 54C = FF
      when "0010101001101" =>  data <= "11111111";  -- 54D = FF
      when "0010101001110" =>  data <= "11111111";  -- 54E = FF
      when "0010101001111" =>  data <= "11111111";  -- 54F = FF
      when "0010101010000" =>  data <= "11111111";  -- 550 = FF
      when "0010101010001" =>  data <= "11111111";  -- 551 = FF
      when "0010101010010" =>  data <= "11111111";  -- 552 = FF
      when "0010101010011" =>  data <= "11111111";  -- 553 = FF
      when "0010101010100" =>  data <= "11111111";  -- 554 = FF
      when "0010101010101" =>  data <= "11111111";  -- 555 = FF
      when "0010101010110" =>  data <= "11111111";  -- 556 = FF
      when "0010101010111" =>  data <= "11111111";  -- 557 = FF
      when "0010101011000" =>  data <= "11111111";  -- 558 = FF
      when "0010101011001" =>  data <= "11111111";  -- 559 = FF
      when "0010101011010" =>  data <= "11111111";  -- 55A = FF
      when "0010101011011" =>  data <= "11111111";  -- 55B = FF
      when "0010101011100" =>  data <= "11111111";  -- 55C = FF
      when "0010101011101" =>  data <= "11111111";  -- 55D = FF
      when "0010101011110" =>  data <= "11111111";  -- 55E = FF
      when "0010101011111" =>  data <= "11111111";  -- 55F = FF
      when "0010101100000" =>  data <= "11111111";  -- 560 = FF
      when "0010101100001" =>  data <= "11111111";  -- 561 = FF
      when "0010101100010" =>  data <= "11111111";  -- 562 = FF
      when "0010101100011" =>  data <= "11111111";  -- 563 = FF
      when "0010101100100" =>  data <= "11111111";  -- 564 = FF
      when "0010101100101" =>  data <= "11111111";  -- 565 = FF
      when "0010101100110" =>  data <= "11111111";  -- 566 = FF
      when "0010101100111" =>  data <= "11111111";  -- 567 = FF
      when "0010101101000" =>  data <= "11111111";  -- 568 = FF
      when "0010101101001" =>  data <= "11111111";  -- 569 = FF
      when "0010101101010" =>  data <= "11111111";  -- 56A = FF
      when "0010101101011" =>  data <= "11111111";  -- 56B = FF
      when "0010101101100" =>  data <= "11111111";  -- 56C = FF
      when "0010101101101" =>  data <= "11111111";  -- 56D = FF
      when "0010101101110" =>  data <= "11111111";  -- 56E = FF
      when "0010101101111" =>  data <= "11111111";  -- 56F = FF
      when "0010101110000" =>  data <= "11111111";  -- 570 = FF
      when "0010101110001" =>  data <= "11111111";  -- 571 = FF
      when "0010101110010" =>  data <= "11111111";  -- 572 = FF
      when "0010101110011" =>  data <= "11111111";  -- 573 = FF
      when "0010101110100" =>  data <= "11111111";  -- 574 = FF
      when "0010101110101" =>  data <= "11111111";  -- 575 = FF
      when "0010101110110" =>  data <= "11111111";  -- 576 = FF
      when "0010101110111" =>  data <= "11111111";  -- 577 = FF
      when "0010101111000" =>  data <= "11111111";  -- 578 = FF
      when "0010101111001" =>  data <= "11111111";  -- 579 = FF
      when "0010101111010" =>  data <= "11111111";  -- 57A = FF
      when "0010101111011" =>  data <= "11111111";  -- 57B = FF
      when "0010101111100" =>  data <= "11111111";  -- 57C = FF
      when "0010101111101" =>  data <= "11111111";  -- 57D = FF
      when "0010101111110" =>  data <= "11111111";  -- 57E = FF
      when "0010101111111" =>  data <= "11111111";  -- 57F = FF
      when "0010110000000" =>  data <= "11111111";  -- 580 = FF
      when "0010110000001" =>  data <= "11111111";  -- 581 = FF
      when "0010110000010" =>  data <= "11111111";  -- 582 = FF
      when "0010110000011" =>  data <= "11111111";  -- 583 = FF
      when "0010110000100" =>  data <= "11111111";  -- 584 = FF
      when "0010110000101" =>  data <= "11111111";  -- 585 = FF
      when "0010110000110" =>  data <= "11111111";  -- 586 = FF
      when "0010110000111" =>  data <= "11111111";  -- 587 = FF
      when "0010110001000" =>  data <= "11111111";  -- 588 = FF
      when "0010110001001" =>  data <= "11111111";  -- 589 = FF
      when "0010110001010" =>  data <= "11111111";  -- 58A = FF
      when "0010110001011" =>  data <= "11111111";  -- 58B = FF
      when "0010110001100" =>  data <= "11111111";  -- 58C = FF
      when "0010110001101" =>  data <= "11111111";  -- 58D = FF
      when "0010110001110" =>  data <= "11111111";  -- 58E = FF
      when "0010110001111" =>  data <= "11111111";  -- 58F = FF
      when "0010110010000" =>  data <= "11111111";  -- 590 = FF
      when "0010110010001" =>  data <= "11111111";  -- 591 = FF
      when "0010110010010" =>  data <= "11111111";  -- 592 = FF
      when "0010110010011" =>  data <= "11111111";  -- 593 = FF
      when "0010110010100" =>  data <= "11111111";  -- 594 = FF
      when "0010110010101" =>  data <= "11111111";  -- 595 = FF
      when "0010110010110" =>  data <= "11111111";  -- 596 = FF
      when "0010110010111" =>  data <= "11111111";  -- 597 = FF
      when "0010110011000" =>  data <= "11111111";  -- 598 = FF
      when "0010110011001" =>  data <= "11111111";  -- 599 = FF
      when "0010110011010" =>  data <= "11111111";  -- 59A = FF
      when "0010110011011" =>  data <= "11111111";  -- 59B = FF
      when "0010110011100" =>  data <= "11111111";  -- 59C = FF
      when "0010110011101" =>  data <= "11111111";  -- 59D = FF
      when "0010110011110" =>  data <= "11111111";  -- 59E = FF
      when "0010110011111" =>  data <= "11111111";  -- 59F = FF
      when "0010110100000" =>  data <= "11111111";  -- 5A0 = FF
      when "0010110100001" =>  data <= "11111111";  -- 5A1 = FF
      when "0010110100010" =>  data <= "11111111";  -- 5A2 = FF
      when "0010110100011" =>  data <= "11111111";  -- 5A3 = FF
      when "0010110100100" =>  data <= "11111111";  -- 5A4 = FF
      when "0010110100101" =>  data <= "11111111";  -- 5A5 = FF
      when "0010110100110" =>  data <= "11111111";  -- 5A6 = FF
      when "0010110100111" =>  data <= "11111111";  -- 5A7 = FF
      when "0010110101000" =>  data <= "11111111";  -- 5A8 = FF
      when "0010110101001" =>  data <= "11111111";  -- 5A9 = FF
      when "0010110101010" =>  data <= "11111111";  -- 5AA = FF
      when "0010110101011" =>  data <= "11111111";  -- 5AB = FF
      when "0010110101100" =>  data <= "11111111";  -- 5AC = FF
      when "0010110101101" =>  data <= "11111111";  -- 5AD = FF
      when "0010110101110" =>  data <= "11111111";  -- 5AE = FF
      when "0010110101111" =>  data <= "11111111";  -- 5AF = FF
      when "0010110110000" =>  data <= "11111111";  -- 5B0 = FF
      when "0010110110001" =>  data <= "11111111";  -- 5B1 = FF
      when "0010110110010" =>  data <= "11111111";  -- 5B2 = FF
      when "0010110110011" =>  data <= "11111111";  -- 5B3 = FF
      when "0010110110100" =>  data <= "11111111";  -- 5B4 = FF
      when "0010110110101" =>  data <= "11111111";  -- 5B5 = FF
      when "0010110110110" =>  data <= "11111111";  -- 5B6 = FF
      when "0010110110111" =>  data <= "11111111";  -- 5B7 = FF
      when "0010110111000" =>  data <= "11111111";  -- 5B8 = FF
      when "0010110111001" =>  data <= "11111111";  -- 5B9 = FF
      when "0010110111010" =>  data <= "11111111";  -- 5BA = FF
      when "0010110111011" =>  data <= "11111111";  -- 5BB = FF
      when "0010110111100" =>  data <= "11111111";  -- 5BC = FF
      when "0010110111101" =>  data <= "11111111";  -- 5BD = FF
      when "0010110111110" =>  data <= "11111111";  -- 5BE = FF
      when "0010110111111" =>  data <= "11111111";  -- 5BF = FF
      when "0010111000000" =>  data <= "11111111";  -- 5C0 = FF
      when "0010111000001" =>  data <= "11111111";  -- 5C1 = FF
      when "0010111000010" =>  data <= "11111111";  -- 5C2 = FF
      when "0010111000011" =>  data <= "11111111";  -- 5C3 = FF
      when "0010111000100" =>  data <= "11111111";  -- 5C4 = FF
      when "0010111000101" =>  data <= "11111111";  -- 5C5 = FF
      when "0010111000110" =>  data <= "11111111";  -- 5C6 = FF
      when "0010111000111" =>  data <= "11111111";  -- 5C7 = FF
      when "0010111001000" =>  data <= "11111111";  -- 5C8 = FF
      when "0010111001001" =>  data <= "11111111";  -- 5C9 = FF
      when "0010111001010" =>  data <= "11111111";  -- 5CA = FF
      when "0010111001011" =>  data <= "11111111";  -- 5CB = FF
      when "0010111001100" =>  data <= "11111111";  -- 5CC = FF
      when "0010111001101" =>  data <= "11111111";  -- 5CD = FF
      when "0010111001110" =>  data <= "11111111";  -- 5CE = FF
      when "0010111001111" =>  data <= "11111111";  -- 5CF = FF
      when "0010111010000" =>  data <= "11111111";  -- 5D0 = FF
      when "0010111010001" =>  data <= "11111111";  -- 5D1 = FF
      when "0010111010010" =>  data <= "11111111";  -- 5D2 = FF
      when "0010111010011" =>  data <= "11111111";  -- 5D3 = FF
      when "0010111010100" =>  data <= "11111111";  -- 5D4 = FF
      when "0010111010101" =>  data <= "11111111";  -- 5D5 = FF
      when "0010111010110" =>  data <= "11111111";  -- 5D6 = FF
      when "0010111010111" =>  data <= "11111111";  -- 5D7 = FF
      when "0010111011000" =>  data <= "11111111";  -- 5D8 = FF
      when "0010111011001" =>  data <= "11111111";  -- 5D9 = FF
      when "0010111011010" =>  data <= "11111111";  -- 5DA = FF
      when "0010111011011" =>  data <= "11111111";  -- 5DB = FF
      when "0010111011100" =>  data <= "11111111";  -- 5DC = FF
      when "0010111011101" =>  data <= "11111111";  -- 5DD = FF
      when "0010111011110" =>  data <= "11111111";  -- 5DE = FF
      when "0010111011111" =>  data <= "11111111";  -- 5DF = FF
      when "0010111100000" =>  data <= "11111111";  -- 5E0 = FF
      when "0010111100001" =>  data <= "11111111";  -- 5E1 = FF
      when "0010111100010" =>  data <= "11111111";  -- 5E2 = FF
      when "0010111100011" =>  data <= "11111111";  -- 5E3 = FF
      when "0010111100100" =>  data <= "11111111";  -- 5E4 = FF
      when "0010111100101" =>  data <= "11111111";  -- 5E5 = FF
      when "0010111100110" =>  data <= "11111111";  -- 5E6 = FF
      when "0010111100111" =>  data <= "11111111";  -- 5E7 = FF
      when "0010111101000" =>  data <= "11111111";  -- 5E8 = FF
      when "0010111101001" =>  data <= "11111111";  -- 5E9 = FF
      when "0010111101010" =>  data <= "11111111";  -- 5EA = FF
      when "0010111101011" =>  data <= "11111111";  -- 5EB = FF
      when "0010111101100" =>  data <= "11111111";  -- 5EC = FF
      when "0010111101101" =>  data <= "11111111";  -- 5ED = FF
      when "0010111101110" =>  data <= "11111111";  -- 5EE = FF
      when "0010111101111" =>  data <= "11111111";  -- 5EF = FF
      when "0010111110000" =>  data <= "11111111";  -- 5F0 = FF
      when "0010111110001" =>  data <= "11111111";  -- 5F1 = FF
      when "0010111110010" =>  data <= "11111111";  -- 5F2 = FF
      when "0010111110011" =>  data <= "11111111";  -- 5F3 = FF
      when "0010111110100" =>  data <= "11111111";  -- 5F4 = FF
      when "0010111110101" =>  data <= "11111111";  -- 5F5 = FF
      when "0010111110110" =>  data <= "11111111";  -- 5F6 = FF
      when "0010111110111" =>  data <= "11111111";  -- 5F7 = FF
      when "0010111111000" =>  data <= "11111111";  -- 5F8 = FF
      when "0010111111001" =>  data <= "11111111";  -- 5F9 = FF
      when "0010111111010" =>  data <= "11111111";  -- 5FA = FF
      when "0010111111011" =>  data <= "11111111";  -- 5FB = FF
      when "0010111111100" =>  data <= "11111111";  -- 5FC = FF
      when "0010111111101" =>  data <= "11111111";  -- 5FD = FF
      when "0010111111110" =>  data <= "11111111";  -- 5FE = FF
      when "0010111111111" =>  data <= "11111111";  -- 5FF = FF
      when "0011000000000" =>  data <= "11111111";  -- 600 = FF
      when "0011000000001" =>  data <= "11111111";  -- 601 = FF
      when "0011000000010" =>  data <= "11111111";  -- 602 = FF
      when "0011000000011" =>  data <= "11111111";  -- 603 = FF
      when "0011000000100" =>  data <= "11111111";  -- 604 = FF
      when "0011000000101" =>  data <= "11111111";  -- 605 = FF
      when "0011000000110" =>  data <= "11111111";  -- 606 = FF
      when "0011000000111" =>  data <= "11111111";  -- 607 = FF
      when "0011000001000" =>  data <= "11111111";  -- 608 = FF
      when "0011000001001" =>  data <= "11111111";  -- 609 = FF
      when "0011000001010" =>  data <= "11111111";  -- 60A = FF
      when "0011000001011" =>  data <= "11111111";  -- 60B = FF
      when "0011000001100" =>  data <= "11111111";  -- 60C = FF
      when "0011000001101" =>  data <= "11111111";  -- 60D = FF
      when "0011000001110" =>  data <= "11111111";  -- 60E = FF
      when "0011000001111" =>  data <= "11111111";  -- 60F = FF
      when "0011000010000" =>  data <= "11111111";  -- 610 = FF
      when "0011000010001" =>  data <= "11111111";  -- 611 = FF
      when "0011000010010" =>  data <= "11111111";  -- 612 = FF
      when "0011000010011" =>  data <= "11111111";  -- 613 = FF
      when "0011000010100" =>  data <= "11111111";  -- 614 = FF
      when "0011000010101" =>  data <= "11111111";  -- 615 = FF
      when "0011000010110" =>  data <= "11111111";  -- 616 = FF
      when "0011000010111" =>  data <= "11111111";  -- 617 = FF
      when "0011000011000" =>  data <= "11111111";  -- 618 = FF
      when "0011000011001" =>  data <= "11111111";  -- 619 = FF
      when "0011000011010" =>  data <= "11111111";  -- 61A = FF
      when "0011000011011" =>  data <= "11111111";  -- 61B = FF
      when "0011000011100" =>  data <= "11111111";  -- 61C = FF
      when "0011000011101" =>  data <= "11111111";  -- 61D = FF
      when "0011000011110" =>  data <= "11111111";  -- 61E = FF
      when "0011000011111" =>  data <= "11111111";  -- 61F = FF
      when "0011000100000" =>  data <= "11111111";  -- 620 = FF
      when "0011000100001" =>  data <= "11111111";  -- 621 = FF
      when "0011000100010" =>  data <= "11111111";  -- 622 = FF
      when "0011000100011" =>  data <= "11111111";  -- 623 = FF
      when "0011000100100" =>  data <= "11111111";  -- 624 = FF
      when "0011000100101" =>  data <= "11111111";  -- 625 = FF
      when "0011000100110" =>  data <= "11111111";  -- 626 = FF
      when "0011000100111" =>  data <= "11111111";  -- 627 = FF
      when "0011000101000" =>  data <= "11111111";  -- 628 = FF
      when "0011000101001" =>  data <= "11111111";  -- 629 = FF
      when "0011000101010" =>  data <= "11111111";  -- 62A = FF
      when "0011000101011" =>  data <= "11111111";  -- 62B = FF
      when "0011000101100" =>  data <= "11111111";  -- 62C = FF
      when "0011000101101" =>  data <= "11111111";  -- 62D = FF
      when "0011000101110" =>  data <= "11111111";  -- 62E = FF
      when "0011000101111" =>  data <= "11111111";  -- 62F = FF
      when "0011000110000" =>  data <= "11111111";  -- 630 = FF
      when "0011000110001" =>  data <= "11111111";  -- 631 = FF
      when "0011000110010" =>  data <= "11111111";  -- 632 = FF
      when "0011000110011" =>  data <= "11111111";  -- 633 = FF
      when "0011000110100" =>  data <= "11111111";  -- 634 = FF
      when "0011000110101" =>  data <= "11111111";  -- 635 = FF
      when "0011000110110" =>  data <= "11111111";  -- 636 = FF
      when "0011000110111" =>  data <= "11111111";  -- 637 = FF
      when "0011000111000" =>  data <= "11111111";  -- 638 = FF
      when "0011000111001" =>  data <= "11111111";  -- 639 = FF
      when "0011000111010" =>  data <= "11111111";  -- 63A = FF
      when "0011000111011" =>  data <= "11111111";  -- 63B = FF
      when "0011000111100" =>  data <= "11111111";  -- 63C = FF
      when "0011000111101" =>  data <= "11111111";  -- 63D = FF
      when "0011000111110" =>  data <= "11111111";  -- 63E = FF
      when "0011000111111" =>  data <= "11111111";  -- 63F = FF
      when "0011001000000" =>  data <= "11111111";  -- 640 = FF
      when "0011001000001" =>  data <= "11111111";  -- 641 = FF
      when "0011001000010" =>  data <= "11111111";  -- 642 = FF
      when "0011001000011" =>  data <= "11111111";  -- 643 = FF
      when "0011001000100" =>  data <= "11111111";  -- 644 = FF
      when "0011001000101" =>  data <= "11111111";  -- 645 = FF
      when "0011001000110" =>  data <= "11111111";  -- 646 = FF
      when "0011001000111" =>  data <= "11111111";  -- 647 = FF
      when "0011001001000" =>  data <= "11111111";  -- 648 = FF
      when "0011001001001" =>  data <= "11111111";  -- 649 = FF
      when "0011001001010" =>  data <= "11111111";  -- 64A = FF
      when "0011001001011" =>  data <= "11111111";  -- 64B = FF
      when "0011001001100" =>  data <= "11111111";  -- 64C = FF
      when "0011001001101" =>  data <= "11111111";  -- 64D = FF
      when "0011001001110" =>  data <= "11111111";  -- 64E = FF
      when "0011001001111" =>  data <= "11111111";  -- 64F = FF
      when "0011001010000" =>  data <= "11111111";  -- 650 = FF
      when "0011001010001" =>  data <= "11111111";  -- 651 = FF
      when "0011001010010" =>  data <= "11111111";  -- 652 = FF
      when "0011001010011" =>  data <= "11111111";  -- 653 = FF
      when "0011001010100" =>  data <= "11111111";  -- 654 = FF
      when "0011001010101" =>  data <= "11111111";  -- 655 = FF
      when "0011001010110" =>  data <= "11111111";  -- 656 = FF
      when "0011001010111" =>  data <= "11111111";  -- 657 = FF
      when "0011001011000" =>  data <= "11111111";  -- 658 = FF
      when "0011001011001" =>  data <= "11111111";  -- 659 = FF
      when "0011001011010" =>  data <= "11111111";  -- 65A = FF
      when "0011001011011" =>  data <= "11111111";  -- 65B = FF
      when "0011001011100" =>  data <= "11111111";  -- 65C = FF
      when "0011001011101" =>  data <= "11111111";  -- 65D = FF
      when "0011001011110" =>  data <= "11111111";  -- 65E = FF
      when "0011001011111" =>  data <= "11111111";  -- 65F = FF
      when "0011001100000" =>  data <= "11111111";  -- 660 = FF
      when "0011001100001" =>  data <= "11111111";  -- 661 = FF
      when "0011001100010" =>  data <= "11111111";  -- 662 = FF
      when "0011001100011" =>  data <= "11111111";  -- 663 = FF
      when "0011001100100" =>  data <= "11111111";  -- 664 = FF
      when "0011001100101" =>  data <= "11111111";  -- 665 = FF
      when "0011001100110" =>  data <= "11111111";  -- 666 = FF
      when "0011001100111" =>  data <= "11111111";  -- 667 = FF
      when "0011001101000" =>  data <= "11111111";  -- 668 = FF
      when "0011001101001" =>  data <= "11111111";  -- 669 = FF
      when "0011001101010" =>  data <= "11111111";  -- 66A = FF
      when "0011001101011" =>  data <= "11111111";  -- 66B = FF
      when "0011001101100" =>  data <= "11111111";  -- 66C = FF
      when "0011001101101" =>  data <= "11111111";  -- 66D = FF
      when "0011001101110" =>  data <= "11111111";  -- 66E = FF
      when "0011001101111" =>  data <= "11111111";  -- 66F = FF
      when "0011001110000" =>  data <= "11111111";  -- 670 = FF
      when "0011001110001" =>  data <= "11111111";  -- 671 = FF
      when "0011001110010" =>  data <= "11111111";  -- 672 = FF
      when "0011001110011" =>  data <= "11111111";  -- 673 = FF
      when "0011001110100" =>  data <= "11111111";  -- 674 = FF
      when "0011001110101" =>  data <= "11111111";  -- 675 = FF
      when "0011001110110" =>  data <= "11111111";  -- 676 = FF
      when "0011001110111" =>  data <= "11111111";  -- 677 = FF
      when "0011001111000" =>  data <= "11111111";  -- 678 = FF
      when "0011001111001" =>  data <= "11111111";  -- 679 = FF
      when "0011001111010" =>  data <= "11111111";  -- 67A = FF
      when "0011001111011" =>  data <= "11111111";  -- 67B = FF
      when "0011001111100" =>  data <= "11111111";  -- 67C = FF
      when "0011001111101" =>  data <= "11111111";  -- 67D = FF
      when "0011001111110" =>  data <= "11111111";  -- 67E = FF
      when "0011001111111" =>  data <= "11111111";  -- 67F = FF
      when "0011010000000" =>  data <= "11111111";  -- 680 = FF
      when "0011010000001" =>  data <= "11111111";  -- 681 = FF
      when "0011010000010" =>  data <= "11111111";  -- 682 = FF
      when "0011010000011" =>  data <= "11111111";  -- 683 = FF
      when "0011010000100" =>  data <= "11111111";  -- 684 = FF
      when "0011010000101" =>  data <= "11111111";  -- 685 = FF
      when "0011010000110" =>  data <= "11111111";  -- 686 = FF
      when "0011010000111" =>  data <= "11111111";  -- 687 = FF
      when "0011010001000" =>  data <= "11111111";  -- 688 = FF
      when "0011010001001" =>  data <= "11111111";  -- 689 = FF
      when "0011010001010" =>  data <= "11111111";  -- 68A = FF
      when "0011010001011" =>  data <= "11111111";  -- 68B = FF
      when "0011010001100" =>  data <= "11111111";  -- 68C = FF
      when "0011010001101" =>  data <= "11111111";  -- 68D = FF
      when "0011010001110" =>  data <= "11111111";  -- 68E = FF
      when "0011010001111" =>  data <= "11111111";  -- 68F = FF
      when "0011010010000" =>  data <= "11111111";  -- 690 = FF
      when "0011010010001" =>  data <= "11111111";  -- 691 = FF
      when "0011010010010" =>  data <= "11111111";  -- 692 = FF
      when "0011010010011" =>  data <= "11111111";  -- 693 = FF
      when "0011010010100" =>  data <= "11111111";  -- 694 = FF
      when "0011010010101" =>  data <= "11111111";  -- 695 = FF
      when "0011010010110" =>  data <= "11111111";  -- 696 = FF
      when "0011010010111" =>  data <= "11111111";  -- 697 = FF
      when "0011010011000" =>  data <= "11111111";  -- 698 = FF
      when "0011010011001" =>  data <= "11111111";  -- 699 = FF
      when "0011010011010" =>  data <= "11111111";  -- 69A = FF
      when "0011010011011" =>  data <= "11111111";  -- 69B = FF
      when "0011010011100" =>  data <= "11111111";  -- 69C = FF
      when "0011010011101" =>  data <= "11111111";  -- 69D = FF
      when "0011010011110" =>  data <= "11111111";  -- 69E = FF
      when "0011010011111" =>  data <= "11111111";  -- 69F = FF
      when "0011010100000" =>  data <= "11111111";  -- 6A0 = FF
      when "0011010100001" =>  data <= "11111111";  -- 6A1 = FF
      when "0011010100010" =>  data <= "11111111";  -- 6A2 = FF
      when "0011010100011" =>  data <= "11111111";  -- 6A3 = FF
      when "0011010100100" =>  data <= "11111111";  -- 6A4 = FF
      when "0011010100101" =>  data <= "11111111";  -- 6A5 = FF
      when "0011010100110" =>  data <= "11111111";  -- 6A6 = FF
      when "0011010100111" =>  data <= "11111111";  -- 6A7 = FF
      when "0011010101000" =>  data <= "11111111";  -- 6A8 = FF
      when "0011010101001" =>  data <= "11111111";  -- 6A9 = FF
      when "0011010101010" =>  data <= "11111111";  -- 6AA = FF
      when "0011010101011" =>  data <= "11111111";  -- 6AB = FF
      when "0011010101100" =>  data <= "11111111";  -- 6AC = FF
      when "0011010101101" =>  data <= "11111111";  -- 6AD = FF
      when "0011010101110" =>  data <= "11111111";  -- 6AE = FF
      when "0011010101111" =>  data <= "11111111";  -- 6AF = FF
      when "0011010110000" =>  data <= "11111111";  -- 6B0 = FF
      when "0011010110001" =>  data <= "11111111";  -- 6B1 = FF
      when "0011010110010" =>  data <= "11111111";  -- 6B2 = FF
      when "0011010110011" =>  data <= "11111111";  -- 6B3 = FF
      when "0011010110100" =>  data <= "11111111";  -- 6B4 = FF
      when "0011010110101" =>  data <= "11111111";  -- 6B5 = FF
      when "0011010110110" =>  data <= "11111111";  -- 6B6 = FF
      when "0011010110111" =>  data <= "11111111";  -- 6B7 = FF
      when "0011010111000" =>  data <= "11111111";  -- 6B8 = FF
      when "0011010111001" =>  data <= "11111111";  -- 6B9 = FF
      when "0011010111010" =>  data <= "11111111";  -- 6BA = FF
      when "0011010111011" =>  data <= "11111111";  -- 6BB = FF
      when "0011010111100" =>  data <= "11111111";  -- 6BC = FF
      when "0011010111101" =>  data <= "11111111";  -- 6BD = FF
      when "0011010111110" =>  data <= "11111111";  -- 6BE = FF
      when "0011010111111" =>  data <= "11111111";  -- 6BF = FF
      when "0011011000000" =>  data <= "11111111";  -- 6C0 = FF
      when "0011011000001" =>  data <= "11111111";  -- 6C1 = FF
      when "0011011000010" =>  data <= "11111111";  -- 6C2 = FF
      when "0011011000011" =>  data <= "11111111";  -- 6C3 = FF
      when "0011011000100" =>  data <= "11111111";  -- 6C4 = FF
      when "0011011000101" =>  data <= "11111111";  -- 6C5 = FF
      when "0011011000110" =>  data <= "11111111";  -- 6C6 = FF
      when "0011011000111" =>  data <= "11111111";  -- 6C7 = FF
      when "0011011001000" =>  data <= "11111111";  -- 6C8 = FF
      when "0011011001001" =>  data <= "11111111";  -- 6C9 = FF
      when "0011011001010" =>  data <= "11111111";  -- 6CA = FF
      when "0011011001011" =>  data <= "11111111";  -- 6CB = FF
      when "0011011001100" =>  data <= "11111111";  -- 6CC = FF
      when "0011011001101" =>  data <= "11111111";  -- 6CD = FF
      when "0011011001110" =>  data <= "11111111";  -- 6CE = FF
      when "0011011001111" =>  data <= "11111111";  -- 6CF = FF
      when "0011011010000" =>  data <= "11111111";  -- 6D0 = FF
      when "0011011010001" =>  data <= "11111111";  -- 6D1 = FF
      when "0011011010010" =>  data <= "11111111";  -- 6D2 = FF
      when "0011011010011" =>  data <= "11111111";  -- 6D3 = FF
      when "0011011010100" =>  data <= "11111111";  -- 6D4 = FF
      when "0011011010101" =>  data <= "11111111";  -- 6D5 = FF
      when "0011011010110" =>  data <= "11111111";  -- 6D6 = FF
      when "0011011010111" =>  data <= "11111111";  -- 6D7 = FF
      when "0011011011000" =>  data <= "11111111";  -- 6D8 = FF
      when "0011011011001" =>  data <= "11111111";  -- 6D9 = FF
      when "0011011011010" =>  data <= "11111111";  -- 6DA = FF
      when "0011011011011" =>  data <= "11111111";  -- 6DB = FF
      when "0011011011100" =>  data <= "11111111";  -- 6DC = FF
      when "0011011011101" =>  data <= "11111111";  -- 6DD = FF
      when "0011011011110" =>  data <= "11111111";  -- 6DE = FF
      when "0011011011111" =>  data <= "11111111";  -- 6DF = FF
      when "0011011100000" =>  data <= "11111111";  -- 6E0 = FF
      when "0011011100001" =>  data <= "11111111";  -- 6E1 = FF
      when "0011011100010" =>  data <= "11111111";  -- 6E2 = FF
      when "0011011100011" =>  data <= "11111111";  -- 6E3 = FF
      when "0011011100100" =>  data <= "11111111";  -- 6E4 = FF
      when "0011011100101" =>  data <= "11111111";  -- 6E5 = FF
      when "0011011100110" =>  data <= "11111111";  -- 6E6 = FF
      when "0011011100111" =>  data <= "11111111";  -- 6E7 = FF
      when "0011011101000" =>  data <= "11111111";  -- 6E8 = FF
      when "0011011101001" =>  data <= "11111111";  -- 6E9 = FF
      when "0011011101010" =>  data <= "11111111";  -- 6EA = FF
      when "0011011101011" =>  data <= "11111111";  -- 6EB = FF
      when "0011011101100" =>  data <= "11111111";  -- 6EC = FF
      when "0011011101101" =>  data <= "11111111";  -- 6ED = FF
      when "0011011101110" =>  data <= "11111111";  -- 6EE = FF
      when "0011011101111" =>  data <= "11111111";  -- 6EF = FF
      when "0011011110000" =>  data <= "11111111";  -- 6F0 = FF
      when "0011011110001" =>  data <= "11111111";  -- 6F1 = FF
      when "0011011110010" =>  data <= "11111111";  -- 6F2 = FF
      when "0011011110011" =>  data <= "11111111";  -- 6F3 = FF
      when "0011011110100" =>  data <= "11111111";  -- 6F4 = FF
      when "0011011110101" =>  data <= "11111111";  -- 6F5 = FF
      when "0011011110110" =>  data <= "11111111";  -- 6F6 = FF
      when "0011011110111" =>  data <= "11111111";  -- 6F7 = FF
      when "0011011111000" =>  data <= "11111111";  -- 6F8 = FF
      when "0011011111001" =>  data <= "11111111";  -- 6F9 = FF
      when "0011011111010" =>  data <= "11111111";  -- 6FA = FF
      when "0011011111011" =>  data <= "11111111";  -- 6FB = FF
      when "0011011111100" =>  data <= "11111111";  -- 6FC = FF
      when "0011011111101" =>  data <= "11111111";  -- 6FD = FF
      when "0011011111110" =>  data <= "11111111";  -- 6FE = FF
      when "0011011111111" =>  data <= "11111111";  -- 6FF = FF
      when "0011100000000" =>  data <= "11111111";  -- 700 = FF
      when "0011100000001" =>  data <= "11111111";  -- 701 = FF
      when "0011100000010" =>  data <= "11111111";  -- 702 = FF
      when "0011100000011" =>  data <= "11111111";  -- 703 = FF
      when "0011100000100" =>  data <= "11111111";  -- 704 = FF
      when "0011100000101" =>  data <= "11111111";  -- 705 = FF
      when "0011100000110" =>  data <= "11111111";  -- 706 = FF
      when "0011100000111" =>  data <= "11111111";  -- 707 = FF
      when "0011100001000" =>  data <= "11111111";  -- 708 = FF
      when "0011100001001" =>  data <= "11111111";  -- 709 = FF
      when "0011100001010" =>  data <= "11111111";  -- 70A = FF
      when "0011100001011" =>  data <= "11111111";  -- 70B = FF
      when "0011100001100" =>  data <= "11111111";  -- 70C = FF
      when "0011100001101" =>  data <= "11111111";  -- 70D = FF
      when "0011100001110" =>  data <= "11111111";  -- 70E = FF
      when "0011100001111" =>  data <= "11111111";  -- 70F = FF
      when "0011100010000" =>  data <= "11111111";  -- 710 = FF
      when "0011100010001" =>  data <= "11111111";  -- 711 = FF
      when "0011100010010" =>  data <= "11111111";  -- 712 = FF
      when "0011100010011" =>  data <= "11111111";  -- 713 = FF
      when "0011100010100" =>  data <= "11111111";  -- 714 = FF
      when "0011100010101" =>  data <= "11111111";  -- 715 = FF
      when "0011100010110" =>  data <= "11111111";  -- 716 = FF
      when "0011100010111" =>  data <= "11111111";  -- 717 = FF
      when "0011100011000" =>  data <= "11111111";  -- 718 = FF
      when "0011100011001" =>  data <= "11111111";  -- 719 = FF
      when "0011100011010" =>  data <= "11111111";  -- 71A = FF
      when "0011100011011" =>  data <= "11111111";  -- 71B = FF
      when "0011100011100" =>  data <= "11111111";  -- 71C = FF
      when "0011100011101" =>  data <= "11111111";  -- 71D = FF
      when "0011100011110" =>  data <= "11111111";  -- 71E = FF
      when "0011100011111" =>  data <= "11111111";  -- 71F = FF
      when "0011100100000" =>  data <= "11111111";  -- 720 = FF
      when "0011100100001" =>  data <= "11111111";  -- 721 = FF
      when "0011100100010" =>  data <= "11111111";  -- 722 = FF
      when "0011100100011" =>  data <= "11111111";  -- 723 = FF
      when "0011100100100" =>  data <= "11111111";  -- 724 = FF
      when "0011100100101" =>  data <= "11111111";  -- 725 = FF
      when "0011100100110" =>  data <= "11111111";  -- 726 = FF
      when "0011100100111" =>  data <= "11111111";  -- 727 = FF
      when "0011100101000" =>  data <= "11111111";  -- 728 = FF
      when "0011100101001" =>  data <= "11111111";  -- 729 = FF
      when "0011100101010" =>  data <= "11111111";  -- 72A = FF
      when "0011100101011" =>  data <= "11111111";  -- 72B = FF
      when "0011100101100" =>  data <= "11111111";  -- 72C = FF
      when "0011100101101" =>  data <= "11111111";  -- 72D = FF
      when "0011100101110" =>  data <= "11111111";  -- 72E = FF
      when "0011100101111" =>  data <= "11111111";  -- 72F = FF
      when "0011100110000" =>  data <= "11111111";  -- 730 = FF
      when "0011100110001" =>  data <= "11111111";  -- 731 = FF
      when "0011100110010" =>  data <= "11111111";  -- 732 = FF
      when "0011100110011" =>  data <= "11111111";  -- 733 = FF
      when "0011100110100" =>  data <= "11111111";  -- 734 = FF
      when "0011100110101" =>  data <= "11111111";  -- 735 = FF
      when "0011100110110" =>  data <= "11111111";  -- 736 = FF
      when "0011100110111" =>  data <= "11111111";  -- 737 = FF
      when "0011100111000" =>  data <= "11111111";  -- 738 = FF
      when "0011100111001" =>  data <= "11111111";  -- 739 = FF
      when "0011100111010" =>  data <= "11111111";  -- 73A = FF
      when "0011100111011" =>  data <= "11111111";  -- 73B = FF
      when "0011100111100" =>  data <= "11111111";  -- 73C = FF
      when "0011100111101" =>  data <= "11111111";  -- 73D = FF
      when "0011100111110" =>  data <= "11111111";  -- 73E = FF
      when "0011100111111" =>  data <= "11111111";  -- 73F = FF
      when "0011101000000" =>  data <= "11111111";  -- 740 = FF
      when "0011101000001" =>  data <= "11111111";  -- 741 = FF
      when "0011101000010" =>  data <= "11111111";  -- 742 = FF
      when "0011101000011" =>  data <= "11111111";  -- 743 = FF
      when "0011101000100" =>  data <= "11111111";  -- 744 = FF
      when "0011101000101" =>  data <= "11111111";  -- 745 = FF
      when "0011101000110" =>  data <= "11111111";  -- 746 = FF
      when "0011101000111" =>  data <= "11111111";  -- 747 = FF
      when "0011101001000" =>  data <= "11111111";  -- 748 = FF
      when "0011101001001" =>  data <= "11111111";  -- 749 = FF
      when "0011101001010" =>  data <= "11111111";  -- 74A = FF
      when "0011101001011" =>  data <= "11111111";  -- 74B = FF
      when "0011101001100" =>  data <= "11111111";  -- 74C = FF
      when "0011101001101" =>  data <= "11111111";  -- 74D = FF
      when "0011101001110" =>  data <= "11111111";  -- 74E = FF
      when "0011101001111" =>  data <= "11111111";  -- 74F = FF
      when "0011101010000" =>  data <= "11111111";  -- 750 = FF
      when "0011101010001" =>  data <= "11111111";  -- 751 = FF
      when "0011101010010" =>  data <= "11111111";  -- 752 = FF
      when "0011101010011" =>  data <= "11111111";  -- 753 = FF
      when "0011101010100" =>  data <= "11111111";  -- 754 = FF
      when "0011101010101" =>  data <= "11111111";  -- 755 = FF
      when "0011101010110" =>  data <= "11111111";  -- 756 = FF
      when "0011101010111" =>  data <= "11111111";  -- 757 = FF
      when "0011101011000" =>  data <= "11111111";  -- 758 = FF
      when "0011101011001" =>  data <= "11111111";  -- 759 = FF
      when "0011101011010" =>  data <= "11111111";  -- 75A = FF
      when "0011101011011" =>  data <= "11111111";  -- 75B = FF
      when "0011101011100" =>  data <= "11111111";  -- 75C = FF
      when "0011101011101" =>  data <= "11111111";  -- 75D = FF
      when "0011101011110" =>  data <= "11111111";  -- 75E = FF
      when "0011101011111" =>  data <= "11111111";  -- 75F = FF
      when "0011101100000" =>  data <= "11111111";  -- 760 = FF
      when "0011101100001" =>  data <= "11111111";  -- 761 = FF
      when "0011101100010" =>  data <= "11111111";  -- 762 = FF
      when "0011101100011" =>  data <= "11111111";  -- 763 = FF
      when "0011101100100" =>  data <= "11111111";  -- 764 = FF
      when "0011101100101" =>  data <= "11111111";  -- 765 = FF
      when "0011101100110" =>  data <= "11111111";  -- 766 = FF
      when "0011101100111" =>  data <= "11111111";  -- 767 = FF
      when "0011101101000" =>  data <= "11111111";  -- 768 = FF
      when "0011101101001" =>  data <= "11111111";  -- 769 = FF
      when "0011101101010" =>  data <= "11111111";  -- 76A = FF
      when "0011101101011" =>  data <= "11111111";  -- 76B = FF
      when "0011101101100" =>  data <= "11111111";  -- 76C = FF
      when "0011101101101" =>  data <= "11111111";  -- 76D = FF
      when "0011101101110" =>  data <= "11111111";  -- 76E = FF
      when "0011101101111" =>  data <= "11111111";  -- 76F = FF
      when "0011101110000" =>  data <= "11111111";  -- 770 = FF
      when "0011101110001" =>  data <= "11111111";  -- 771 = FF
      when "0011101110010" =>  data <= "11111111";  -- 772 = FF
      when "0011101110011" =>  data <= "11111111";  -- 773 = FF
      when "0011101110100" =>  data <= "11111111";  -- 774 = FF
      when "0011101110101" =>  data <= "11111111";  -- 775 = FF
      when "0011101110110" =>  data <= "11111111";  -- 776 = FF
      when "0011101110111" =>  data <= "11111111";  -- 777 = FF
      when "0011101111000" =>  data <= "11111111";  -- 778 = FF
      when "0011101111001" =>  data <= "11111111";  -- 779 = FF
      when "0011101111010" =>  data <= "11111111";  -- 77A = FF
      when "0011101111011" =>  data <= "11111111";  -- 77B = FF
      when "0011101111100" =>  data <= "11111111";  -- 77C = FF
      when "0011101111101" =>  data <= "11111111";  -- 77D = FF
      when "0011101111110" =>  data <= "11111111";  -- 77E = FF
      when "0011101111111" =>  data <= "11111111";  -- 77F = FF
      when "0011110000000" =>  data <= "11111111";  -- 780 = FF
      when "0011110000001" =>  data <= "11111111";  -- 781 = FF
      when "0011110000010" =>  data <= "11111111";  -- 782 = FF
      when "0011110000011" =>  data <= "11111111";  -- 783 = FF
      when "0011110000100" =>  data <= "11111111";  -- 784 = FF
      when "0011110000101" =>  data <= "11111111";  -- 785 = FF
      when "0011110000110" =>  data <= "11111111";  -- 786 = FF
      when "0011110000111" =>  data <= "11111111";  -- 787 = FF
      when "0011110001000" =>  data <= "11111111";  -- 788 = FF
      when "0011110001001" =>  data <= "11111111";  -- 789 = FF
      when "0011110001010" =>  data <= "11111111";  -- 78A = FF
      when "0011110001011" =>  data <= "11111111";  -- 78B = FF
      when "0011110001100" =>  data <= "11111111";  -- 78C = FF
      when "0011110001101" =>  data <= "11111111";  -- 78D = FF
      when "0011110001110" =>  data <= "11111111";  -- 78E = FF
      when "0011110001111" =>  data <= "11111111";  -- 78F = FF
      when "0011110010000" =>  data <= "11111111";  -- 790 = FF
      when "0011110010001" =>  data <= "11111111";  -- 791 = FF
      when "0011110010010" =>  data <= "11111111";  -- 792 = FF
      when "0011110010011" =>  data <= "11111111";  -- 793 = FF
      when "0011110010100" =>  data <= "11111111";  -- 794 = FF
      when "0011110010101" =>  data <= "11111111";  -- 795 = FF
      when "0011110010110" =>  data <= "11111111";  -- 796 = FF
      when "0011110010111" =>  data <= "11111111";  -- 797 = FF
      when "0011110011000" =>  data <= "11111111";  -- 798 = FF
      when "0011110011001" =>  data <= "11111111";  -- 799 = FF
      when "0011110011010" =>  data <= "11111111";  -- 79A = FF
      when "0011110011011" =>  data <= "11111111";  -- 79B = FF
      when "0011110011100" =>  data <= "11111111";  -- 79C = FF
      when "0011110011101" =>  data <= "11111111";  -- 79D = FF
      when "0011110011110" =>  data <= "11111111";  -- 79E = FF
      when "0011110011111" =>  data <= "11111111";  -- 79F = FF
      when "0011110100000" =>  data <= "11111111";  -- 7A0 = FF
      when "0011110100001" =>  data <= "11111111";  -- 7A1 = FF
      when "0011110100010" =>  data <= "11111111";  -- 7A2 = FF
      when "0011110100011" =>  data <= "11111111";  -- 7A3 = FF
      when "0011110100100" =>  data <= "11111111";  -- 7A4 = FF
      when "0011110100101" =>  data <= "11111111";  -- 7A5 = FF
      when "0011110100110" =>  data <= "11111111";  -- 7A6 = FF
      when "0011110100111" =>  data <= "11111111";  -- 7A7 = FF
      when "0011110101000" =>  data <= "11111111";  -- 7A8 = FF
      when "0011110101001" =>  data <= "11111111";  -- 7A9 = FF
      when "0011110101010" =>  data <= "11111111";  -- 7AA = FF
      when "0011110101011" =>  data <= "11111111";  -- 7AB = FF
      when "0011110101100" =>  data <= "11111111";  -- 7AC = FF
      when "0011110101101" =>  data <= "11111111";  -- 7AD = FF
      when "0011110101110" =>  data <= "11111111";  -- 7AE = FF
      when "0011110101111" =>  data <= "11111111";  -- 7AF = FF
      when "0011110110000" =>  data <= "11111111";  -- 7B0 = FF
      when "0011110110001" =>  data <= "11111111";  -- 7B1 = FF
      when "0011110110010" =>  data <= "11111111";  -- 7B2 = FF
      when "0011110110011" =>  data <= "11111111";  -- 7B3 = FF
      when "0011110110100" =>  data <= "11111111";  -- 7B4 = FF
      when "0011110110101" =>  data <= "11111111";  -- 7B5 = FF
      when "0011110110110" =>  data <= "11111111";  -- 7B6 = FF
      when "0011110110111" =>  data <= "11111111";  -- 7B7 = FF
      when "0011110111000" =>  data <= "11111111";  -- 7B8 = FF
      when "0011110111001" =>  data <= "11111111";  -- 7B9 = FF
      when "0011110111010" =>  data <= "11111111";  -- 7BA = FF
      when "0011110111011" =>  data <= "11111111";  -- 7BB = FF
      when "0011110111100" =>  data <= "11111111";  -- 7BC = FF
      when "0011110111101" =>  data <= "11111111";  -- 7BD = FF
      when "0011110111110" =>  data <= "11111111";  -- 7BE = FF
      when "0011110111111" =>  data <= "11111111";  -- 7BF = FF
      when "0011111000000" =>  data <= "11111111";  -- 7C0 = FF
      when "0011111000001" =>  data <= "11111111";  -- 7C1 = FF
      when "0011111000010" =>  data <= "11111111";  -- 7C2 = FF
      when "0011111000011" =>  data <= "11111111";  -- 7C3 = FF
      when "0011111000100" =>  data <= "11111111";  -- 7C4 = FF
      when "0011111000101" =>  data <= "11111111";  -- 7C5 = FF
      when "0011111000110" =>  data <= "11111111";  -- 7C6 = FF
      when "0011111000111" =>  data <= "11111111";  -- 7C7 = FF
      when "0011111001000" =>  data <= "11111111";  -- 7C8 = FF
      when "0011111001001" =>  data <= "11111111";  -- 7C9 = FF
      when "0011111001010" =>  data <= "11111111";  -- 7CA = FF
      when "0011111001011" =>  data <= "11111111";  -- 7CB = FF
      when "0011111001100" =>  data <= "11111111";  -- 7CC = FF
      when "0011111001101" =>  data <= "11111111";  -- 7CD = FF
      when "0011111001110" =>  data <= "11111111";  -- 7CE = FF
      when "0011111001111" =>  data <= "11111111";  -- 7CF = FF
      when "0011111010000" =>  data <= "11111111";  -- 7D0 = FF
      when "0011111010001" =>  data <= "11111111";  -- 7D1 = FF
      when "0011111010010" =>  data <= "11111111";  -- 7D2 = FF
      when "0011111010011" =>  data <= "11111111";  -- 7D3 = FF
      when "0011111010100" =>  data <= "11111111";  -- 7D4 = FF
      when "0011111010101" =>  data <= "11111111";  -- 7D5 = FF
      when "0011111010110" =>  data <= "11111111";  -- 7D6 = FF
      when "0011111010111" =>  data <= "11111111";  -- 7D7 = FF
      when "0011111011000" =>  data <= "11111111";  -- 7D8 = FF
      when "0011111011001" =>  data <= "11111111";  -- 7D9 = FF
      when "0011111011010" =>  data <= "11111111";  -- 7DA = FF
      when "0011111011011" =>  data <= "11111111";  -- 7DB = FF
      when "0011111011100" =>  data <= "11111111";  -- 7DC = FF
      when "0011111011101" =>  data <= "11111111";  -- 7DD = FF
      when "0011111011110" =>  data <= "11111111";  -- 7DE = FF
      when "0011111011111" =>  data <= "11111111";  -- 7DF = FF
      when "0011111100000" =>  data <= "11111111";  -- 7E0 = FF
      when "0011111100001" =>  data <= "11111111";  -- 7E1 = FF
      when "0011111100010" =>  data <= "11111111";  -- 7E2 = FF
      when "0011111100011" =>  data <= "11111111";  -- 7E3 = FF
      when "0011111100100" =>  data <= "11111111";  -- 7E4 = FF
      when "0011111100101" =>  data <= "11111111";  -- 7E5 = FF
      when "0011111100110" =>  data <= "11111111";  -- 7E6 = FF
      when "0011111100111" =>  data <= "11111111";  -- 7E7 = FF
      when "0011111101000" =>  data <= "11111111";  -- 7E8 = FF
      when "0011111101001" =>  data <= "11111111";  -- 7E9 = FF
      when "0011111101010" =>  data <= "11111111";  -- 7EA = FF
      when "0011111101011" =>  data <= "11111111";  -- 7EB = FF
      when "0011111101100" =>  data <= "11111111";  -- 7EC = FF
      when "0011111101101" =>  data <= "11111111";  -- 7ED = FF
      when "0011111101110" =>  data <= "11111111";  -- 7EE = FF
      when "0011111101111" =>  data <= "11111111";  -- 7EF = FF
      when "0011111110000" =>  data <= "11111111";  -- 7F0 = FF
      when "0011111110001" =>  data <= "11111111";  -- 7F1 = FF
      when "0011111110010" =>  data <= "11111111";  -- 7F2 = FF
      when "0011111110011" =>  data <= "11111111";  -- 7F3 = FF
      when "0011111110100" =>  data <= "11111111";  -- 7F4 = FF
      when "0011111110101" =>  data <= "11111111";  -- 7F5 = FF
      when "0011111110110" =>  data <= "11111111";  -- 7F6 = FF
      when "0011111110111" =>  data <= "11111111";  -- 7F7 = FF
      when "0011111111000" =>  data <= "11111111";  -- 7F8 = FF
      when "0011111111001" =>  data <= "11111111";  -- 7F9 = FF
      when "0011111111010" =>  data <= "11111111";  -- 7FA = FF
      when "0011111111011" =>  data <= "11111111";  -- 7FB = FF
      when "0011111111100" =>  data <= "11111111";  -- 7FC = FF
      when "0011111111101" =>  data <= "11111111";  -- 7FD = FF
      when "0011111111110" =>  data <= "11111111";  -- 7FE = FF
      when "0011111111111" =>  data <= "11111111";  -- 7FF = FF
      when "0100000000000" =>  data <= "11111111";  -- 800 = FF
      when "0100000000001" =>  data <= "11111111";  -- 801 = FF
      when "0100000000010" =>  data <= "11111111";  -- 802 = FF
      when "0100000000011" =>  data <= "11111111";  -- 803 = FF
      when "0100000000100" =>  data <= "11111111";  -- 804 = FF
      when "0100000000101" =>  data <= "11111111";  -- 805 = FF
      when "0100000000110" =>  data <= "11111111";  -- 806 = FF
      when "0100000000111" =>  data <= "11111111";  -- 807 = FF
      when "0100000001000" =>  data <= "11111111";  -- 808 = FF
      when "0100000001001" =>  data <= "11111111";  -- 809 = FF
      when "0100000001010" =>  data <= "11111111";  -- 80A = FF
      when "0100000001011" =>  data <= "11111111";  -- 80B = FF
      when "0100000001100" =>  data <= "11111111";  -- 80C = FF
      when "0100000001101" =>  data <= "11111111";  -- 80D = FF
      when "0100000001110" =>  data <= "11111111";  -- 80E = FF
      when "0100000001111" =>  data <= "11111111";  -- 80F = FF
      when "0100000010000" =>  data <= "11111111";  -- 810 = FF
      when "0100000010001" =>  data <= "11111111";  -- 811 = FF
      when "0100000010010" =>  data <= "11111111";  -- 812 = FF
      when "0100000010011" =>  data <= "11111111";  -- 813 = FF
      when "0100000010100" =>  data <= "11111111";  -- 814 = FF
      when "0100000010101" =>  data <= "11111111";  -- 815 = FF
      when "0100000010110" =>  data <= "11111111";  -- 816 = FF
      when "0100000010111" =>  data <= "11111111";  -- 817 = FF
      when "0100000011000" =>  data <= "11111111";  -- 818 = FF
      when "0100000011001" =>  data <= "11111111";  -- 819 = FF
      when "0100000011010" =>  data <= "11111111";  -- 81A = FF
      when "0100000011011" =>  data <= "11111111";  -- 81B = FF
      when "0100000011100" =>  data <= "11111111";  -- 81C = FF
      when "0100000011101" =>  data <= "11111111";  -- 81D = FF
      when "0100000011110" =>  data <= "11111111";  -- 81E = FF
      when "0100000011111" =>  data <= "11111111";  -- 81F = FF
      when "0100000100000" =>  data <= "11111111";  -- 820 = FF
      when "0100000100001" =>  data <= "11111111";  -- 821 = FF
      when "0100000100010" =>  data <= "11111111";  -- 822 = FF
      when "0100000100011" =>  data <= "11111111";  -- 823 = FF
      when "0100000100100" =>  data <= "11111111";  -- 824 = FF
      when "0100000100101" =>  data <= "11111111";  -- 825 = FF
      when "0100000100110" =>  data <= "11111111";  -- 826 = FF
      when "0100000100111" =>  data <= "11111111";  -- 827 = FF
      when "0100000101000" =>  data <= "11111111";  -- 828 = FF
      when "0100000101001" =>  data <= "11111111";  -- 829 = FF
      when "0100000101010" =>  data <= "11111111";  -- 82A = FF
      when "0100000101011" =>  data <= "11111111";  -- 82B = FF
      when "0100000101100" =>  data <= "11111111";  -- 82C = FF
      when "0100000101101" =>  data <= "11111111";  -- 82D = FF
      when "0100000101110" =>  data <= "11111111";  -- 82E = FF
      when "0100000101111" =>  data <= "11111111";  -- 82F = FF
      when "0100000110000" =>  data <= "11111111";  -- 830 = FF
      when "0100000110001" =>  data <= "11111111";  -- 831 = FF
      when "0100000110010" =>  data <= "11111111";  -- 832 = FF
      when "0100000110011" =>  data <= "11111111";  -- 833 = FF
      when "0100000110100" =>  data <= "11111111";  -- 834 = FF
      when "0100000110101" =>  data <= "11111111";  -- 835 = FF
      when "0100000110110" =>  data <= "11111111";  -- 836 = FF
      when "0100000110111" =>  data <= "11111111";  -- 837 = FF
      when "0100000111000" =>  data <= "11111111";  -- 838 = FF
      when "0100000111001" =>  data <= "11111111";  -- 839 = FF
      when "0100000111010" =>  data <= "11111111";  -- 83A = FF
      when "0100000111011" =>  data <= "11111111";  -- 83B = FF
      when "0100000111100" =>  data <= "11111111";  -- 83C = FF
      when "0100000111101" =>  data <= "11111111";  -- 83D = FF
      when "0100000111110" =>  data <= "11111111";  -- 83E = FF
      when "0100000111111" =>  data <= "11111111";  -- 83F = FF
      when "0100001000000" =>  data <= "11111111";  -- 840 = FF
      when "0100001000001" =>  data <= "11111111";  -- 841 = FF
      when "0100001000010" =>  data <= "11111111";  -- 842 = FF
      when "0100001000011" =>  data <= "11111111";  -- 843 = FF
      when "0100001000100" =>  data <= "11111111";  -- 844 = FF
      when "0100001000101" =>  data <= "11111111";  -- 845 = FF
      when "0100001000110" =>  data <= "11111111";  -- 846 = FF
      when "0100001000111" =>  data <= "11111111";  -- 847 = FF
      when "0100001001000" =>  data <= "11111111";  -- 848 = FF
      when "0100001001001" =>  data <= "11111111";  -- 849 = FF
      when "0100001001010" =>  data <= "11111111";  -- 84A = FF
      when "0100001001011" =>  data <= "11111111";  -- 84B = FF
      when "0100001001100" =>  data <= "11111111";  -- 84C = FF
      when "0100001001101" =>  data <= "11111111";  -- 84D = FF
      when "0100001001110" =>  data <= "11111111";  -- 84E = FF
      when "0100001001111" =>  data <= "11111111";  -- 84F = FF
      when "0100001010000" =>  data <= "11111111";  -- 850 = FF
      when "0100001010001" =>  data <= "11111111";  -- 851 = FF
      when "0100001010010" =>  data <= "11111111";  -- 852 = FF
      when "0100001010011" =>  data <= "11111111";  -- 853 = FF
      when "0100001010100" =>  data <= "11111111";  -- 854 = FF
      when "0100001010101" =>  data <= "11111111";  -- 855 = FF
      when "0100001010110" =>  data <= "11111111";  -- 856 = FF
      when "0100001010111" =>  data <= "11111111";  -- 857 = FF
      when "0100001011000" =>  data <= "11111111";  -- 858 = FF
      when "0100001011001" =>  data <= "11111111";  -- 859 = FF
      when "0100001011010" =>  data <= "11111111";  -- 85A = FF
      when "0100001011011" =>  data <= "11111111";  -- 85B = FF
      when "0100001011100" =>  data <= "11111111";  -- 85C = FF
      when "0100001011101" =>  data <= "11111111";  -- 85D = FF
      when "0100001011110" =>  data <= "11111111";  -- 85E = FF
      when "0100001011111" =>  data <= "11111111";  -- 85F = FF
      when "0100001100000" =>  data <= "11111111";  -- 860 = FF
      when "0100001100001" =>  data <= "11111111";  -- 861 = FF
      when "0100001100010" =>  data <= "11111111";  -- 862 = FF
      when "0100001100011" =>  data <= "11111111";  -- 863 = FF
      when "0100001100100" =>  data <= "11111111";  -- 864 = FF
      when "0100001100101" =>  data <= "11111111";  -- 865 = FF
      when "0100001100110" =>  data <= "11111111";  -- 866 = FF
      when "0100001100111" =>  data <= "11111111";  -- 867 = FF
      when "0100001101000" =>  data <= "11111111";  -- 868 = FF
      when "0100001101001" =>  data <= "11111111";  -- 869 = FF
      when "0100001101010" =>  data <= "11111111";  -- 86A = FF
      when "0100001101011" =>  data <= "11111111";  -- 86B = FF
      when "0100001101100" =>  data <= "11111111";  -- 86C = FF
      when "0100001101101" =>  data <= "11111111";  -- 86D = FF
      when "0100001101110" =>  data <= "11111111";  -- 86E = FF
      when "0100001101111" =>  data <= "11111111";  -- 86F = FF
      when "0100001110000" =>  data <= "11111111";  -- 870 = FF
      when "0100001110001" =>  data <= "11111111";  -- 871 = FF
      when "0100001110010" =>  data <= "11111111";  -- 872 = FF
      when "0100001110011" =>  data <= "11111111";  -- 873 = FF
      when "0100001110100" =>  data <= "11111111";  -- 874 = FF
      when "0100001110101" =>  data <= "11111111";  -- 875 = FF
      when "0100001110110" =>  data <= "11111111";  -- 876 = FF
      when "0100001110111" =>  data <= "11111111";  -- 877 = FF
      when "0100001111000" =>  data <= "11111111";  -- 878 = FF
      when "0100001111001" =>  data <= "11111111";  -- 879 = FF
      when "0100001111010" =>  data <= "11111111";  -- 87A = FF
      when "0100001111011" =>  data <= "11111111";  -- 87B = FF
      when "0100001111100" =>  data <= "11111111";  -- 87C = FF
      when "0100001111101" =>  data <= "11111111";  -- 87D = FF
      when "0100001111110" =>  data <= "11111111";  -- 87E = FF
      when "0100001111111" =>  data <= "11111111";  -- 87F = FF
      when "0100010000000" =>  data <= "11111111";  -- 880 = FF
      when "0100010000001" =>  data <= "11111111";  -- 881 = FF
      when "0100010000010" =>  data <= "11111111";  -- 882 = FF
      when "0100010000011" =>  data <= "11111111";  -- 883 = FF
      when "0100010000100" =>  data <= "11111111";  -- 884 = FF
      when "0100010000101" =>  data <= "11111111";  -- 885 = FF
      when "0100010000110" =>  data <= "11111111";  -- 886 = FF
      when "0100010000111" =>  data <= "11111111";  -- 887 = FF
      when "0100010001000" =>  data <= "11111111";  -- 888 = FF
      when "0100010001001" =>  data <= "11111111";  -- 889 = FF
      when "0100010001010" =>  data <= "11111111";  -- 88A = FF
      when "0100010001011" =>  data <= "11111111";  -- 88B = FF
      when "0100010001100" =>  data <= "11111111";  -- 88C = FF
      when "0100010001101" =>  data <= "11111111";  -- 88D = FF
      when "0100010001110" =>  data <= "11111111";  -- 88E = FF
      when "0100010001111" =>  data <= "11111111";  -- 88F = FF
      when "0100010010000" =>  data <= "11111111";  -- 890 = FF
      when "0100010010001" =>  data <= "11111111";  -- 891 = FF
      when "0100010010010" =>  data <= "11111111";  -- 892 = FF
      when "0100010010011" =>  data <= "11111111";  -- 893 = FF
      when "0100010010100" =>  data <= "11111111";  -- 894 = FF
      when "0100010010101" =>  data <= "11111111";  -- 895 = FF
      when "0100010010110" =>  data <= "11111111";  -- 896 = FF
      when "0100010010111" =>  data <= "11111111";  -- 897 = FF
      when "0100010011000" =>  data <= "11111111";  -- 898 = FF
      when "0100010011001" =>  data <= "11111111";  -- 899 = FF
      when "0100010011010" =>  data <= "11111111";  -- 89A = FF
      when "0100010011011" =>  data <= "11111111";  -- 89B = FF
      when "0100010011100" =>  data <= "11111111";  -- 89C = FF
      when "0100010011101" =>  data <= "11111111";  -- 89D = FF
      when "0100010011110" =>  data <= "11111111";  -- 89E = FF
      when "0100010011111" =>  data <= "11111111";  -- 89F = FF
      when "0100010100000" =>  data <= "11111111";  -- 8A0 = FF
      when "0100010100001" =>  data <= "11111111";  -- 8A1 = FF
      when "0100010100010" =>  data <= "11111111";  -- 8A2 = FF
      when "0100010100011" =>  data <= "11111111";  -- 8A3 = FF
      when "0100010100100" =>  data <= "11111111";  -- 8A4 = FF
      when "0100010100101" =>  data <= "11111111";  -- 8A5 = FF
      when "0100010100110" =>  data <= "11111111";  -- 8A6 = FF
      when "0100010100111" =>  data <= "11111111";  -- 8A7 = FF
      when "0100010101000" =>  data <= "11111111";  -- 8A8 = FF
      when "0100010101001" =>  data <= "11111111";  -- 8A9 = FF
      when "0100010101010" =>  data <= "11111111";  -- 8AA = FF
      when "0100010101011" =>  data <= "11111111";  -- 8AB = FF
      when "0100010101100" =>  data <= "11111111";  -- 8AC = FF
      when "0100010101101" =>  data <= "11111111";  -- 8AD = FF
      when "0100010101110" =>  data <= "11111111";  -- 8AE = FF
      when "0100010101111" =>  data <= "11111111";  -- 8AF = FF
      when "0100010110000" =>  data <= "11111111";  -- 8B0 = FF
      when "0100010110001" =>  data <= "11111111";  -- 8B1 = FF
      when "0100010110010" =>  data <= "11111111";  -- 8B2 = FF
      when "0100010110011" =>  data <= "11111111";  -- 8B3 = FF
      when "0100010110100" =>  data <= "11111111";  -- 8B4 = FF
      when "0100010110101" =>  data <= "11111111";  -- 8B5 = FF
      when "0100010110110" =>  data <= "11111111";  -- 8B6 = FF
      when "0100010110111" =>  data <= "11111111";  -- 8B7 = FF
      when "0100010111000" =>  data <= "11111111";  -- 8B8 = FF
      when "0100010111001" =>  data <= "11111111";  -- 8B9 = FF
      when "0100010111010" =>  data <= "11111111";  -- 8BA = FF
      when "0100010111011" =>  data <= "11111111";  -- 8BB = FF
      when "0100010111100" =>  data <= "11111111";  -- 8BC = FF
      when "0100010111101" =>  data <= "11111111";  -- 8BD = FF
      when "0100010111110" =>  data <= "11111111";  -- 8BE = FF
      when "0100010111111" =>  data <= "11111111";  -- 8BF = FF
      when "0100011000000" =>  data <= "11111111";  -- 8C0 = FF
      when "0100011000001" =>  data <= "11111111";  -- 8C1 = FF
      when "0100011000010" =>  data <= "11111111";  -- 8C2 = FF
      when "0100011000011" =>  data <= "11111111";  -- 8C3 = FF
      when "0100011000100" =>  data <= "11111111";  -- 8C4 = FF
      when "0100011000101" =>  data <= "11111111";  -- 8C5 = FF
      when "0100011000110" =>  data <= "11111111";  -- 8C6 = FF
      when "0100011000111" =>  data <= "11111111";  -- 8C7 = FF
      when "0100011001000" =>  data <= "11111111";  -- 8C8 = FF
      when "0100011001001" =>  data <= "11111111";  -- 8C9 = FF
      when "0100011001010" =>  data <= "11111111";  -- 8CA = FF
      when "0100011001011" =>  data <= "11111111";  -- 8CB = FF
      when "0100011001100" =>  data <= "11111111";  -- 8CC = FF
      when "0100011001101" =>  data <= "11111111";  -- 8CD = FF
      when "0100011001110" =>  data <= "11111111";  -- 8CE = FF
      when "0100011001111" =>  data <= "11111111";  -- 8CF = FF
      when "0100011010000" =>  data <= "11111111";  -- 8D0 = FF
      when "0100011010001" =>  data <= "11111111";  -- 8D1 = FF
      when "0100011010010" =>  data <= "11111111";  -- 8D2 = FF
      when "0100011010011" =>  data <= "11111111";  -- 8D3 = FF
      when "0100011010100" =>  data <= "11111111";  -- 8D4 = FF
      when "0100011010101" =>  data <= "11111111";  -- 8D5 = FF
      when "0100011010110" =>  data <= "11111111";  -- 8D6 = FF
      when "0100011010111" =>  data <= "11111111";  -- 8D7 = FF
      when "0100011011000" =>  data <= "11111111";  -- 8D8 = FF
      when "0100011011001" =>  data <= "11111111";  -- 8D9 = FF
      when "0100011011010" =>  data <= "11111111";  -- 8DA = FF
      when "0100011011011" =>  data <= "11111111";  -- 8DB = FF
      when "0100011011100" =>  data <= "11111111";  -- 8DC = FF
      when "0100011011101" =>  data <= "11111111";  -- 8DD = FF
      when "0100011011110" =>  data <= "11111111";  -- 8DE = FF
      when "0100011011111" =>  data <= "11111111";  -- 8DF = FF
      when "0100011100000" =>  data <= "11111111";  -- 8E0 = FF
      when "0100011100001" =>  data <= "11111111";  -- 8E1 = FF
      when "0100011100010" =>  data <= "11111111";  -- 8E2 = FF
      when "0100011100011" =>  data <= "11111111";  -- 8E3 = FF
      when "0100011100100" =>  data <= "11111111";  -- 8E4 = FF
      when "0100011100101" =>  data <= "11111111";  -- 8E5 = FF
      when "0100011100110" =>  data <= "11111111";  -- 8E6 = FF
      when "0100011100111" =>  data <= "11111111";  -- 8E7 = FF
      when "0100011101000" =>  data <= "11111111";  -- 8E8 = FF
      when "0100011101001" =>  data <= "11111111";  -- 8E9 = FF
      when "0100011101010" =>  data <= "11111111";  -- 8EA = FF
      when "0100011101011" =>  data <= "11111111";  -- 8EB = FF
      when "0100011101100" =>  data <= "11111111";  -- 8EC = FF
      when "0100011101101" =>  data <= "11111111";  -- 8ED = FF
      when "0100011101110" =>  data <= "11111111";  -- 8EE = FF
      when "0100011101111" =>  data <= "11111111";  -- 8EF = FF
      when "0100011110000" =>  data <= "11111111";  -- 8F0 = FF
      when "0100011110001" =>  data <= "11111111";  -- 8F1 = FF
      when "0100011110010" =>  data <= "11111111";  -- 8F2 = FF
      when "0100011110011" =>  data <= "11111111";  -- 8F3 = FF
      when "0100011110100" =>  data <= "11111111";  -- 8F4 = FF
      when "0100011110101" =>  data <= "11111111";  -- 8F5 = FF
      when "0100011110110" =>  data <= "11111111";  -- 8F6 = FF
      when "0100011110111" =>  data <= "11111111";  -- 8F7 = FF
      when "0100011111000" =>  data <= "11111111";  -- 8F8 = FF
      when "0100011111001" =>  data <= "11111111";  -- 8F9 = FF
      when "0100011111010" =>  data <= "11111111";  -- 8FA = FF
      when "0100011111011" =>  data <= "11111111";  -- 8FB = FF
      when "0100011111100" =>  data <= "11111111";  -- 8FC = FF
      when "0100011111101" =>  data <= "11111111";  -- 8FD = FF
      when "0100011111110" =>  data <= "11111111";  -- 8FE = FF
      when "0100011111111" =>  data <= "11111111";  -- 8FF = FF
      when "0100100000000" =>  data <= "11111111";  -- 900 = FF
      when "0100100000001" =>  data <= "11111111";  -- 901 = FF
      when "0100100000010" =>  data <= "11111111";  -- 902 = FF
      when "0100100000011" =>  data <= "11111111";  -- 903 = FF
      when "0100100000100" =>  data <= "11111111";  -- 904 = FF
      when "0100100000101" =>  data <= "11111111";  -- 905 = FF
      when "0100100000110" =>  data <= "11111111";  -- 906 = FF
      when "0100100000111" =>  data <= "11111111";  -- 907 = FF
      when "0100100001000" =>  data <= "11111111";  -- 908 = FF
      when "0100100001001" =>  data <= "11111111";  -- 909 = FF
      when "0100100001010" =>  data <= "11111111";  -- 90A = FF
      when "0100100001011" =>  data <= "11111111";  -- 90B = FF
      when "0100100001100" =>  data <= "11111111";  -- 90C = FF
      when "0100100001101" =>  data <= "11111111";  -- 90D = FF
      when "0100100001110" =>  data <= "11111111";  -- 90E = FF
      when "0100100001111" =>  data <= "11111111";  -- 90F = FF
      when "0100100010000" =>  data <= "11111111";  -- 910 = FF
      when "0100100010001" =>  data <= "11111111";  -- 911 = FF
      when "0100100010010" =>  data <= "11111111";  -- 912 = FF
      when "0100100010011" =>  data <= "11111111";  -- 913 = FF
      when "0100100010100" =>  data <= "11111111";  -- 914 = FF
      when "0100100010101" =>  data <= "11111111";  -- 915 = FF
      when "0100100010110" =>  data <= "11111111";  -- 916 = FF
      when "0100100010111" =>  data <= "11111111";  -- 917 = FF
      when "0100100011000" =>  data <= "11111111";  -- 918 = FF
      when "0100100011001" =>  data <= "11111111";  -- 919 = FF
      when "0100100011010" =>  data <= "11111111";  -- 91A = FF
      when "0100100011011" =>  data <= "11111111";  -- 91B = FF
      when "0100100011100" =>  data <= "11111111";  -- 91C = FF
      when "0100100011101" =>  data <= "11111111";  -- 91D = FF
      when "0100100011110" =>  data <= "11111111";  -- 91E = FF
      when "0100100011111" =>  data <= "11111111";  -- 91F = FF
      when "0100100100000" =>  data <= "11111111";  -- 920 = FF
      when "0100100100001" =>  data <= "11111111";  -- 921 = FF
      when "0100100100010" =>  data <= "11111111";  -- 922 = FF
      when "0100100100011" =>  data <= "11111111";  -- 923 = FF
      when "0100100100100" =>  data <= "11111111";  -- 924 = FF
      when "0100100100101" =>  data <= "11111111";  -- 925 = FF
      when "0100100100110" =>  data <= "11111111";  -- 926 = FF
      when "0100100100111" =>  data <= "11111111";  -- 927 = FF
      when "0100100101000" =>  data <= "11111111";  -- 928 = FF
      when "0100100101001" =>  data <= "11111111";  -- 929 = FF
      when "0100100101010" =>  data <= "11111111";  -- 92A = FF
      when "0100100101011" =>  data <= "11111111";  -- 92B = FF
      when "0100100101100" =>  data <= "11111111";  -- 92C = FF
      when "0100100101101" =>  data <= "11111111";  -- 92D = FF
      when "0100100101110" =>  data <= "11111111";  -- 92E = FF
      when "0100100101111" =>  data <= "11111111";  -- 92F = FF
      when "0100100110000" =>  data <= "11111111";  -- 930 = FF
      when "0100100110001" =>  data <= "11111111";  -- 931 = FF
      when "0100100110010" =>  data <= "11111111";  -- 932 = FF
      when "0100100110011" =>  data <= "11111111";  -- 933 = FF
      when "0100100110100" =>  data <= "11111111";  -- 934 = FF
      when "0100100110101" =>  data <= "11111111";  -- 935 = FF
      when "0100100110110" =>  data <= "11111111";  -- 936 = FF
      when "0100100110111" =>  data <= "11111111";  -- 937 = FF
      when "0100100111000" =>  data <= "11111111";  -- 938 = FF
      when "0100100111001" =>  data <= "11111111";  -- 939 = FF
      when "0100100111010" =>  data <= "11111111";  -- 93A = FF
      when "0100100111011" =>  data <= "11111111";  -- 93B = FF
      when "0100100111100" =>  data <= "11111111";  -- 93C = FF
      when "0100100111101" =>  data <= "11111111";  -- 93D = FF
      when "0100100111110" =>  data <= "11111111";  -- 93E = FF
      when "0100100111111" =>  data <= "11111111";  -- 93F = FF
      when "0100101000000" =>  data <= "11111111";  -- 940 = FF
      when "0100101000001" =>  data <= "11111111";  -- 941 = FF
      when "0100101000010" =>  data <= "11111111";  -- 942 = FF
      when "0100101000011" =>  data <= "11111111";  -- 943 = FF
      when "0100101000100" =>  data <= "11111111";  -- 944 = FF
      when "0100101000101" =>  data <= "11111111";  -- 945 = FF
      when "0100101000110" =>  data <= "11111111";  -- 946 = FF
      when "0100101000111" =>  data <= "11111111";  -- 947 = FF
      when "0100101001000" =>  data <= "11111111";  -- 948 = FF
      when "0100101001001" =>  data <= "11111111";  -- 949 = FF
      when "0100101001010" =>  data <= "11111111";  -- 94A = FF
      when "0100101001011" =>  data <= "11111111";  -- 94B = FF
      when "0100101001100" =>  data <= "11111111";  -- 94C = FF
      when "0100101001101" =>  data <= "11111111";  -- 94D = FF
      when "0100101001110" =>  data <= "11111111";  -- 94E = FF
      when "0100101001111" =>  data <= "11111111";  -- 94F = FF
      when "0100101010000" =>  data <= "11111111";  -- 950 = FF
      when "0100101010001" =>  data <= "11111111";  -- 951 = FF
      when "0100101010010" =>  data <= "11111111";  -- 952 = FF
      when "0100101010011" =>  data <= "11111111";  -- 953 = FF
      when "0100101010100" =>  data <= "11111111";  -- 954 = FF
      when "0100101010101" =>  data <= "11111111";  -- 955 = FF
      when "0100101010110" =>  data <= "11111111";  -- 956 = FF
      when "0100101010111" =>  data <= "11111111";  -- 957 = FF
      when "0100101011000" =>  data <= "11111111";  -- 958 = FF
      when "0100101011001" =>  data <= "11111111";  -- 959 = FF
      when "0100101011010" =>  data <= "11111111";  -- 95A = FF
      when "0100101011011" =>  data <= "11111111";  -- 95B = FF
      when "0100101011100" =>  data <= "11111111";  -- 95C = FF
      when "0100101011101" =>  data <= "11111111";  -- 95D = FF
      when "0100101011110" =>  data <= "11111111";  -- 95E = FF
      when "0100101011111" =>  data <= "11111111";  -- 95F = FF
      when "0100101100000" =>  data <= "11111111";  -- 960 = FF
      when "0100101100001" =>  data <= "11111111";  -- 961 = FF
      when "0100101100010" =>  data <= "11111111";  -- 962 = FF
      when "0100101100011" =>  data <= "11111111";  -- 963 = FF
      when "0100101100100" =>  data <= "11111111";  -- 964 = FF
      when "0100101100101" =>  data <= "11111111";  -- 965 = FF
      when "0100101100110" =>  data <= "11111111";  -- 966 = FF
      when "0100101100111" =>  data <= "11111111";  -- 967 = FF
      when "0100101101000" =>  data <= "11111111";  -- 968 = FF
      when "0100101101001" =>  data <= "11111111";  -- 969 = FF
      when "0100101101010" =>  data <= "11111111";  -- 96A = FF
      when "0100101101011" =>  data <= "11111111";  -- 96B = FF
      when "0100101101100" =>  data <= "11111111";  -- 96C = FF
      when "0100101101101" =>  data <= "11111111";  -- 96D = FF
      when "0100101101110" =>  data <= "11111111";  -- 96E = FF
      when "0100101101111" =>  data <= "11111111";  -- 96F = FF
      when "0100101110000" =>  data <= "11111111";  -- 970 = FF
      when "0100101110001" =>  data <= "11111111";  -- 971 = FF
      when "0100101110010" =>  data <= "11111111";  -- 972 = FF
      when "0100101110011" =>  data <= "11111111";  -- 973 = FF
      when "0100101110100" =>  data <= "11111111";  -- 974 = FF
      when "0100101110101" =>  data <= "11111111";  -- 975 = FF
      when "0100101110110" =>  data <= "11111111";  -- 976 = FF
      when "0100101110111" =>  data <= "11111111";  -- 977 = FF
      when "0100101111000" =>  data <= "11111111";  -- 978 = FF
      when "0100101111001" =>  data <= "11111111";  -- 979 = FF
      when "0100101111010" =>  data <= "11111111";  -- 97A = FF
      when "0100101111011" =>  data <= "11111111";  -- 97B = FF
      when "0100101111100" =>  data <= "11111111";  -- 97C = FF
      when "0100101111101" =>  data <= "11111111";  -- 97D = FF
      when "0100101111110" =>  data <= "11111111";  -- 97E = FF
      when "0100101111111" =>  data <= "11111111";  -- 97F = FF
      when "0100110000000" =>  data <= "11111111";  -- 980 = FF
      when "0100110000001" =>  data <= "11111111";  -- 981 = FF
      when "0100110000010" =>  data <= "11111111";  -- 982 = FF
      when "0100110000011" =>  data <= "11111111";  -- 983 = FF
      when "0100110000100" =>  data <= "11111111";  -- 984 = FF
      when "0100110000101" =>  data <= "11111111";  -- 985 = FF
      when "0100110000110" =>  data <= "11111111";  -- 986 = FF
      when "0100110000111" =>  data <= "11111111";  -- 987 = FF
      when "0100110001000" =>  data <= "11111111";  -- 988 = FF
      when "0100110001001" =>  data <= "11111111";  -- 989 = FF
      when "0100110001010" =>  data <= "11111111";  -- 98A = FF
      when "0100110001011" =>  data <= "11111111";  -- 98B = FF
      when "0100110001100" =>  data <= "11111111";  -- 98C = FF
      when "0100110001101" =>  data <= "11111111";  -- 98D = FF
      when "0100110001110" =>  data <= "11111111";  -- 98E = FF
      when "0100110001111" =>  data <= "11111111";  -- 98F = FF
      when "0100110010000" =>  data <= "11111111";  -- 990 = FF
      when "0100110010001" =>  data <= "11111111";  -- 991 = FF
      when "0100110010010" =>  data <= "11111111";  -- 992 = FF
      when "0100110010011" =>  data <= "11111111";  -- 993 = FF
      when "0100110010100" =>  data <= "11111111";  -- 994 = FF
      when "0100110010101" =>  data <= "11111111";  -- 995 = FF
      when "0100110010110" =>  data <= "11111111";  -- 996 = FF
      when "0100110010111" =>  data <= "11111111";  -- 997 = FF
      when "0100110011000" =>  data <= "11111111";  -- 998 = FF
      when "0100110011001" =>  data <= "11111111";  -- 999 = FF
      when "0100110011010" =>  data <= "11111111";  -- 99A = FF
      when "0100110011011" =>  data <= "11111111";  -- 99B = FF
      when "0100110011100" =>  data <= "11111111";  -- 99C = FF
      when "0100110011101" =>  data <= "11111111";  -- 99D = FF
      when "0100110011110" =>  data <= "11111111";  -- 99E = FF
      when "0100110011111" =>  data <= "11111111";  -- 99F = FF
      when "0100110100000" =>  data <= "11111111";  -- 9A0 = FF
      when "0100110100001" =>  data <= "11111111";  -- 9A1 = FF
      when "0100110100010" =>  data <= "11111111";  -- 9A2 = FF
      when "0100110100011" =>  data <= "11111111";  -- 9A3 = FF
      when "0100110100100" =>  data <= "11111111";  -- 9A4 = FF
      when "0100110100101" =>  data <= "11111111";  -- 9A5 = FF
      when "0100110100110" =>  data <= "11111111";  -- 9A6 = FF
      when "0100110100111" =>  data <= "11111111";  -- 9A7 = FF
      when "0100110101000" =>  data <= "11111111";  -- 9A8 = FF
      when "0100110101001" =>  data <= "11111111";  -- 9A9 = FF
      when "0100110101010" =>  data <= "11111111";  -- 9AA = FF
      when "0100110101011" =>  data <= "11111111";  -- 9AB = FF
      when "0100110101100" =>  data <= "11111111";  -- 9AC = FF
      when "0100110101101" =>  data <= "11111111";  -- 9AD = FF
      when "0100110101110" =>  data <= "11111111";  -- 9AE = FF
      when "0100110101111" =>  data <= "11111111";  -- 9AF = FF
      when "0100110110000" =>  data <= "11111111";  -- 9B0 = FF
      when "0100110110001" =>  data <= "11111111";  -- 9B1 = FF
      when "0100110110010" =>  data <= "11111111";  -- 9B2 = FF
      when "0100110110011" =>  data <= "11111111";  -- 9B3 = FF
      when "0100110110100" =>  data <= "11111111";  -- 9B4 = FF
      when "0100110110101" =>  data <= "11111111";  -- 9B5 = FF
      when "0100110110110" =>  data <= "11111111";  -- 9B6 = FF
      when "0100110110111" =>  data <= "11111111";  -- 9B7 = FF
      when "0100110111000" =>  data <= "11111111";  -- 9B8 = FF
      when "0100110111001" =>  data <= "11111111";  -- 9B9 = FF
      when "0100110111010" =>  data <= "11111111";  -- 9BA = FF
      when "0100110111011" =>  data <= "11111111";  -- 9BB = FF
      when "0100110111100" =>  data <= "11111111";  -- 9BC = FF
      when "0100110111101" =>  data <= "11111111";  -- 9BD = FF
      when "0100110111110" =>  data <= "11111111";  -- 9BE = FF
      when "0100110111111" =>  data <= "11111111";  -- 9BF = FF
      when "0100111000000" =>  data <= "11111111";  -- 9C0 = FF
      when "0100111000001" =>  data <= "11111111";  -- 9C1 = FF
      when "0100111000010" =>  data <= "11111111";  -- 9C2 = FF
      when "0100111000011" =>  data <= "11111111";  -- 9C3 = FF
      when "0100111000100" =>  data <= "11111111";  -- 9C4 = FF
      when "0100111000101" =>  data <= "11111111";  -- 9C5 = FF
      when "0100111000110" =>  data <= "11111111";  -- 9C6 = FF
      when "0100111000111" =>  data <= "11111111";  -- 9C7 = FF
      when "0100111001000" =>  data <= "11111111";  -- 9C8 = FF
      when "0100111001001" =>  data <= "11111111";  -- 9C9 = FF
      when "0100111001010" =>  data <= "11111111";  -- 9CA = FF
      when "0100111001011" =>  data <= "11111111";  -- 9CB = FF
      when "0100111001100" =>  data <= "11111111";  -- 9CC = FF
      when "0100111001101" =>  data <= "11111111";  -- 9CD = FF
      when "0100111001110" =>  data <= "11111111";  -- 9CE = FF
      when "0100111001111" =>  data <= "11111111";  -- 9CF = FF
      when "0100111010000" =>  data <= "11111111";  -- 9D0 = FF
      when "0100111010001" =>  data <= "11111111";  -- 9D1 = FF
      when "0100111010010" =>  data <= "11111111";  -- 9D2 = FF
      when "0100111010011" =>  data <= "11111111";  -- 9D3 = FF
      when "0100111010100" =>  data <= "11111111";  -- 9D4 = FF
      when "0100111010101" =>  data <= "11111111";  -- 9D5 = FF
      when "0100111010110" =>  data <= "11111111";  -- 9D6 = FF
      when "0100111010111" =>  data <= "11111111";  -- 9D7 = FF
      when "0100111011000" =>  data <= "11111111";  -- 9D8 = FF
      when "0100111011001" =>  data <= "11111111";  -- 9D9 = FF
      when "0100111011010" =>  data <= "11111111";  -- 9DA = FF
      when "0100111011011" =>  data <= "11111111";  -- 9DB = FF
      when "0100111011100" =>  data <= "11111111";  -- 9DC = FF
      when "0100111011101" =>  data <= "11111111";  -- 9DD = FF
      when "0100111011110" =>  data <= "11111111";  -- 9DE = FF
      when "0100111011111" =>  data <= "11111111";  -- 9DF = FF
      when "0100111100000" =>  data <= "11111111";  -- 9E0 = FF
      when "0100111100001" =>  data <= "11111111";  -- 9E1 = FF
      when "0100111100010" =>  data <= "11111111";  -- 9E2 = FF
      when "0100111100011" =>  data <= "11111111";  -- 9E3 = FF
      when "0100111100100" =>  data <= "11111111";  -- 9E4 = FF
      when "0100111100101" =>  data <= "11111111";  -- 9E5 = FF
      when "0100111100110" =>  data <= "11111111";  -- 9E6 = FF
      when "0100111100111" =>  data <= "11111111";  -- 9E7 = FF
      when "0100111101000" =>  data <= "11111111";  -- 9E8 = FF
      when "0100111101001" =>  data <= "11111111";  -- 9E9 = FF
      when "0100111101010" =>  data <= "11111111";  -- 9EA = FF
      when "0100111101011" =>  data <= "11111111";  -- 9EB = FF
      when "0100111101100" =>  data <= "11111111";  -- 9EC = FF
      when "0100111101101" =>  data <= "11111111";  -- 9ED = FF
      when "0100111101110" =>  data <= "11111111";  -- 9EE = FF
      when "0100111101111" =>  data <= "11111111";  -- 9EF = FF
      when "0100111110000" =>  data <= "11111111";  -- 9F0 = FF
      when "0100111110001" =>  data <= "11111111";  -- 9F1 = FF
      when "0100111110010" =>  data <= "11111111";  -- 9F2 = FF
      when "0100111110011" =>  data <= "11111111";  -- 9F3 = FF
      when "0100111110100" =>  data <= "11111111";  -- 9F4 = FF
      when "0100111110101" =>  data <= "11111111";  -- 9F5 = FF
      when "0100111110110" =>  data <= "11111111";  -- 9F6 = FF
      when "0100111110111" =>  data <= "11111111";  -- 9F7 = FF
      when "0100111111000" =>  data <= "11111111";  -- 9F8 = FF
      when "0100111111001" =>  data <= "11111111";  -- 9F9 = FF
      when "0100111111010" =>  data <= "11111111";  -- 9FA = FF
      when "0100111111011" =>  data <= "11111111";  -- 9FB = FF
      when "0100111111100" =>  data <= "11111111";  -- 9FC = FF
      when "0100111111101" =>  data <= "11111111";  -- 9FD = FF
      when "0100111111110" =>  data <= "11111111";  -- 9FE = FF
      when "0100111111111" =>  data <= "11111111";  -- 9FF = FF
      when "0101000000000" =>  data <= "11111111";  -- A00 = FF
      when "0101000000001" =>  data <= "11111111";  -- A01 = FF
      when "0101000000010" =>  data <= "11111111";  -- A02 = FF
      when "0101000000011" =>  data <= "11111111";  -- A03 = FF
      when "0101000000100" =>  data <= "11111111";  -- A04 = FF
      when "0101000000101" =>  data <= "11111111";  -- A05 = FF
      when "0101000000110" =>  data <= "11111111";  -- A06 = FF
      when "0101000000111" =>  data <= "11111111";  -- A07 = FF
      when "0101000001000" =>  data <= "11111111";  -- A08 = FF
      when "0101000001001" =>  data <= "11111111";  -- A09 = FF
      when "0101000001010" =>  data <= "11111111";  -- A0A = FF
      when "0101000001011" =>  data <= "11111111";  -- A0B = FF
      when "0101000001100" =>  data <= "11111111";  -- A0C = FF
      when "0101000001101" =>  data <= "11111111";  -- A0D = FF
      when "0101000001110" =>  data <= "11111111";  -- A0E = FF
      when "0101000001111" =>  data <= "11111111";  -- A0F = FF
      when "0101000010000" =>  data <= "11111111";  -- A10 = FF
      when "0101000010001" =>  data <= "11111111";  -- A11 = FF
      when "0101000010010" =>  data <= "11111111";  -- A12 = FF
      when "0101000010011" =>  data <= "11111111";  -- A13 = FF
      when "0101000010100" =>  data <= "11111111";  -- A14 = FF
      when "0101000010101" =>  data <= "11111111";  -- A15 = FF
      when "0101000010110" =>  data <= "11111111";  -- A16 = FF
      when "0101000010111" =>  data <= "11111111";  -- A17 = FF
      when "0101000011000" =>  data <= "11111111";  -- A18 = FF
      when "0101000011001" =>  data <= "11111111";  -- A19 = FF
      when "0101000011010" =>  data <= "11111111";  -- A1A = FF
      when "0101000011011" =>  data <= "11111111";  -- A1B = FF
      when "0101000011100" =>  data <= "11111111";  -- A1C = FF
      when "0101000011101" =>  data <= "11111111";  -- A1D = FF
      when "0101000011110" =>  data <= "11111111";  -- A1E = FF
      when "0101000011111" =>  data <= "11111111";  -- A1F = FF
      when "0101000100000" =>  data <= "11111111";  -- A20 = FF
      when "0101000100001" =>  data <= "11111111";  -- A21 = FF
      when "0101000100010" =>  data <= "11111111";  -- A22 = FF
      when "0101000100011" =>  data <= "11111111";  -- A23 = FF
      when "0101000100100" =>  data <= "11111111";  -- A24 = FF
      when "0101000100101" =>  data <= "11111111";  -- A25 = FF
      when "0101000100110" =>  data <= "11111111";  -- A26 = FF
      when "0101000100111" =>  data <= "11111111";  -- A27 = FF
      when "0101000101000" =>  data <= "11111111";  -- A28 = FF
      when "0101000101001" =>  data <= "11111111";  -- A29 = FF
      when "0101000101010" =>  data <= "11111111";  -- A2A = FF
      when "0101000101011" =>  data <= "11111111";  -- A2B = FF
      when "0101000101100" =>  data <= "11111111";  -- A2C = FF
      when "0101000101101" =>  data <= "11111111";  -- A2D = FF
      when "0101000101110" =>  data <= "11111111";  -- A2E = FF
      when "0101000101111" =>  data <= "11111111";  -- A2F = FF
      when "0101000110000" =>  data <= "11111111";  -- A30 = FF
      when "0101000110001" =>  data <= "11111111";  -- A31 = FF
      when "0101000110010" =>  data <= "11111111";  -- A32 = FF
      when "0101000110011" =>  data <= "11111111";  -- A33 = FF
      when "0101000110100" =>  data <= "11111111";  -- A34 = FF
      when "0101000110101" =>  data <= "11111111";  -- A35 = FF
      when "0101000110110" =>  data <= "11111111";  -- A36 = FF
      when "0101000110111" =>  data <= "11111111";  -- A37 = FF
      when "0101000111000" =>  data <= "11111111";  -- A38 = FF
      when "0101000111001" =>  data <= "11111111";  -- A39 = FF
      when "0101000111010" =>  data <= "11111111";  -- A3A = FF
      when "0101000111011" =>  data <= "11111111";  -- A3B = FF
      when "0101000111100" =>  data <= "11111111";  -- A3C = FF
      when "0101000111101" =>  data <= "11111111";  -- A3D = FF
      when "0101000111110" =>  data <= "11111111";  -- A3E = FF
      when "0101000111111" =>  data <= "11111111";  -- A3F = FF
      when "0101001000000" =>  data <= "11111111";  -- A40 = FF
      when "0101001000001" =>  data <= "11111111";  -- A41 = FF
      when "0101001000010" =>  data <= "11111111";  -- A42 = FF
      when "0101001000011" =>  data <= "11111111";  -- A43 = FF
      when "0101001000100" =>  data <= "11111111";  -- A44 = FF
      when "0101001000101" =>  data <= "11111111";  -- A45 = FF
      when "0101001000110" =>  data <= "11111111";  -- A46 = FF
      when "0101001000111" =>  data <= "11111111";  -- A47 = FF
      when "0101001001000" =>  data <= "11111111";  -- A48 = FF
      when "0101001001001" =>  data <= "11111111";  -- A49 = FF
      when "0101001001010" =>  data <= "11111111";  -- A4A = FF
      when "0101001001011" =>  data <= "11111111";  -- A4B = FF
      when "0101001001100" =>  data <= "11111111";  -- A4C = FF
      when "0101001001101" =>  data <= "11111111";  -- A4D = FF
      when "0101001001110" =>  data <= "11111111";  -- A4E = FF
      when "0101001001111" =>  data <= "11111111";  -- A4F = FF
      when "0101001010000" =>  data <= "11111111";  -- A50 = FF
      when "0101001010001" =>  data <= "11111111";  -- A51 = FF
      when "0101001010010" =>  data <= "11111111";  -- A52 = FF
      when "0101001010011" =>  data <= "11111111";  -- A53 = FF
      when "0101001010100" =>  data <= "11111111";  -- A54 = FF
      when "0101001010101" =>  data <= "11111111";  -- A55 = FF
      when "0101001010110" =>  data <= "11111111";  -- A56 = FF
      when "0101001010111" =>  data <= "11111111";  -- A57 = FF
      when "0101001011000" =>  data <= "11111111";  -- A58 = FF
      when "0101001011001" =>  data <= "11111111";  -- A59 = FF
      when "0101001011010" =>  data <= "11111111";  -- A5A = FF
      when "0101001011011" =>  data <= "11111111";  -- A5B = FF
      when "0101001011100" =>  data <= "11111111";  -- A5C = FF
      when "0101001011101" =>  data <= "11111111";  -- A5D = FF
      when "0101001011110" =>  data <= "11111111";  -- A5E = FF
      when "0101001011111" =>  data <= "11111111";  -- A5F = FF
      when "0101001100000" =>  data <= "11111111";  -- A60 = FF
      when "0101001100001" =>  data <= "11111111";  -- A61 = FF
      when "0101001100010" =>  data <= "11111111";  -- A62 = FF
      when "0101001100011" =>  data <= "11111111";  -- A63 = FF
      when "0101001100100" =>  data <= "11111111";  -- A64 = FF
      when "0101001100101" =>  data <= "11111111";  -- A65 = FF
      when "0101001100110" =>  data <= "11111111";  -- A66 = FF
      when "0101001100111" =>  data <= "11111111";  -- A67 = FF
      when "0101001101000" =>  data <= "11111111";  -- A68 = FF
      when "0101001101001" =>  data <= "11111111";  -- A69 = FF
      when "0101001101010" =>  data <= "11111111";  -- A6A = FF
      when "0101001101011" =>  data <= "11111111";  -- A6B = FF
      when "0101001101100" =>  data <= "11111111";  -- A6C = FF
      when "0101001101101" =>  data <= "11111111";  -- A6D = FF
      when "0101001101110" =>  data <= "11111111";  -- A6E = FF
      when "0101001101111" =>  data <= "11111111";  -- A6F = FF
      when "0101001110000" =>  data <= "11111111";  -- A70 = FF
      when "0101001110001" =>  data <= "11111111";  -- A71 = FF
      when "0101001110010" =>  data <= "11111111";  -- A72 = FF
      when "0101001110011" =>  data <= "11111111";  -- A73 = FF
      when "0101001110100" =>  data <= "11111111";  -- A74 = FF
      when "0101001110101" =>  data <= "11111111";  -- A75 = FF
      when "0101001110110" =>  data <= "11111111";  -- A76 = FF
      when "0101001110111" =>  data <= "11111111";  -- A77 = FF
      when "0101001111000" =>  data <= "11111111";  -- A78 = FF
      when "0101001111001" =>  data <= "11111111";  -- A79 = FF
      when "0101001111010" =>  data <= "11111111";  -- A7A = FF
      when "0101001111011" =>  data <= "11111111";  -- A7B = FF
      when "0101001111100" =>  data <= "11111111";  -- A7C = FF
      when "0101001111101" =>  data <= "11111111";  -- A7D = FF
      when "0101001111110" =>  data <= "11111111";  -- A7E = FF
      when "0101001111111" =>  data <= "11111111";  -- A7F = FF
      when "0101010000000" =>  data <= "11111111";  -- A80 = FF
      when "0101010000001" =>  data <= "11111111";  -- A81 = FF
      when "0101010000010" =>  data <= "11111111";  -- A82 = FF
      when "0101010000011" =>  data <= "11111111";  -- A83 = FF
      when "0101010000100" =>  data <= "11111111";  -- A84 = FF
      when "0101010000101" =>  data <= "11111111";  -- A85 = FF
      when "0101010000110" =>  data <= "11111111";  -- A86 = FF
      when "0101010000111" =>  data <= "11111111";  -- A87 = FF
      when "0101010001000" =>  data <= "11111111";  -- A88 = FF
      when "0101010001001" =>  data <= "11111111";  -- A89 = FF
      when "0101010001010" =>  data <= "11111111";  -- A8A = FF
      when "0101010001011" =>  data <= "11111111";  -- A8B = FF
      when "0101010001100" =>  data <= "11111111";  -- A8C = FF
      when "0101010001101" =>  data <= "11111111";  -- A8D = FF
      when "0101010001110" =>  data <= "11111111";  -- A8E = FF
      when "0101010001111" =>  data <= "11111111";  -- A8F = FF
      when "0101010010000" =>  data <= "11111111";  -- A90 = FF
      when "0101010010001" =>  data <= "11111111";  -- A91 = FF
      when "0101010010010" =>  data <= "11111111";  -- A92 = FF
      when "0101010010011" =>  data <= "11111111";  -- A93 = FF
      when "0101010010100" =>  data <= "11111111";  -- A94 = FF
      when "0101010010101" =>  data <= "11111111";  -- A95 = FF
      when "0101010010110" =>  data <= "11111111";  -- A96 = FF
      when "0101010010111" =>  data <= "11111111";  -- A97 = FF
      when "0101010011000" =>  data <= "11111111";  -- A98 = FF
      when "0101010011001" =>  data <= "11111111";  -- A99 = FF
      when "0101010011010" =>  data <= "11111111";  -- A9A = FF
      when "0101010011011" =>  data <= "11111111";  -- A9B = FF
      when "0101010011100" =>  data <= "11111111";  -- A9C = FF
      when "0101010011101" =>  data <= "11111111";  -- A9D = FF
      when "0101010011110" =>  data <= "11111111";  -- A9E = FF
      when "0101010011111" =>  data <= "11111111";  -- A9F = FF
      when "0101010100000" =>  data <= "11111111";  -- AA0 = FF
      when "0101010100001" =>  data <= "11111111";  -- AA1 = FF
      when "0101010100010" =>  data <= "11111111";  -- AA2 = FF
      when "0101010100011" =>  data <= "11111111";  -- AA3 = FF
      when "0101010100100" =>  data <= "11111111";  -- AA4 = FF
      when "0101010100101" =>  data <= "11111111";  -- AA5 = FF
      when "0101010100110" =>  data <= "11111111";  -- AA6 = FF
      when "0101010100111" =>  data <= "11111111";  -- AA7 = FF
      when "0101010101000" =>  data <= "11111111";  -- AA8 = FF
      when "0101010101001" =>  data <= "11111111";  -- AA9 = FF
      when "0101010101010" =>  data <= "11111111";  -- AAA = FF
      when "0101010101011" =>  data <= "11111111";  -- AAB = FF
      when "0101010101100" =>  data <= "11111111";  -- AAC = FF
      when "0101010101101" =>  data <= "11111111";  -- AAD = FF
      when "0101010101110" =>  data <= "11111111";  -- AAE = FF
      when "0101010101111" =>  data <= "11111111";  -- AAF = FF
      when "0101010110000" =>  data <= "11111111";  -- AB0 = FF
      when "0101010110001" =>  data <= "11111111";  -- AB1 = FF
      when "0101010110010" =>  data <= "11111111";  -- AB2 = FF
      when "0101010110011" =>  data <= "11111111";  -- AB3 = FF
      when "0101010110100" =>  data <= "11111111";  -- AB4 = FF
      when "0101010110101" =>  data <= "11111111";  -- AB5 = FF
      when "0101010110110" =>  data <= "11111111";  -- AB6 = FF
      when "0101010110111" =>  data <= "11111111";  -- AB7 = FF
      when "0101010111000" =>  data <= "11111111";  -- AB8 = FF
      when "0101010111001" =>  data <= "11111111";  -- AB9 = FF
      when "0101010111010" =>  data <= "11111111";  -- ABA = FF
      when "0101010111011" =>  data <= "11111111";  -- ABB = FF
      when "0101010111100" =>  data <= "11111111";  -- ABC = FF
      when "0101010111101" =>  data <= "11111111";  -- ABD = FF
      when "0101010111110" =>  data <= "11111111";  -- ABE = FF
      when "0101010111111" =>  data <= "11111111";  -- ABF = FF
      when "0101011000000" =>  data <= "11111111";  -- AC0 = FF
      when "0101011000001" =>  data <= "11111111";  -- AC1 = FF
      when "0101011000010" =>  data <= "11111111";  -- AC2 = FF
      when "0101011000011" =>  data <= "11111111";  -- AC3 = FF
      when "0101011000100" =>  data <= "11111111";  -- AC4 = FF
      when "0101011000101" =>  data <= "11111111";  -- AC5 = FF
      when "0101011000110" =>  data <= "11111111";  -- AC6 = FF
      when "0101011000111" =>  data <= "11111111";  -- AC7 = FF
      when "0101011001000" =>  data <= "11111111";  -- AC8 = FF
      when "0101011001001" =>  data <= "11111111";  -- AC9 = FF
      when "0101011001010" =>  data <= "11111111";  -- ACA = FF
      when "0101011001011" =>  data <= "11111111";  -- ACB = FF
      when "0101011001100" =>  data <= "11111111";  -- ACC = FF
      when "0101011001101" =>  data <= "11111111";  -- ACD = FF
      when "0101011001110" =>  data <= "11111111";  -- ACE = FF
      when "0101011001111" =>  data <= "11111111";  -- ACF = FF
      when "0101011010000" =>  data <= "11111111";  -- AD0 = FF
      when "0101011010001" =>  data <= "11111111";  -- AD1 = FF
      when "0101011010010" =>  data <= "11111111";  -- AD2 = FF
      when "0101011010011" =>  data <= "11111111";  -- AD3 = FF
      when "0101011010100" =>  data <= "11111111";  -- AD4 = FF
      when "0101011010101" =>  data <= "11111111";  -- AD5 = FF
      when "0101011010110" =>  data <= "11111111";  -- AD6 = FF
      when "0101011010111" =>  data <= "11111111";  -- AD7 = FF
      when "0101011011000" =>  data <= "11111111";  -- AD8 = FF
      when "0101011011001" =>  data <= "11111111";  -- AD9 = FF
      when "0101011011010" =>  data <= "11111111";  -- ADA = FF
      when "0101011011011" =>  data <= "11111111";  -- ADB = FF
      when "0101011011100" =>  data <= "11111111";  -- ADC = FF
      when "0101011011101" =>  data <= "11111111";  -- ADD = FF
      when "0101011011110" =>  data <= "11111111";  -- ADE = FF
      when "0101011011111" =>  data <= "11111111";  -- ADF = FF
      when "0101011100000" =>  data <= "11111111";  -- AE0 = FF
      when "0101011100001" =>  data <= "11111111";  -- AE1 = FF
      when "0101011100010" =>  data <= "11111111";  -- AE2 = FF
      when "0101011100011" =>  data <= "11111111";  -- AE3 = FF
      when "0101011100100" =>  data <= "11111111";  -- AE4 = FF
      when "0101011100101" =>  data <= "11111111";  -- AE5 = FF
      when "0101011100110" =>  data <= "11111111";  -- AE6 = FF
      when "0101011100111" =>  data <= "11111111";  -- AE7 = FF
      when "0101011101000" =>  data <= "11111111";  -- AE8 = FF
      when "0101011101001" =>  data <= "11111111";  -- AE9 = FF
      when "0101011101010" =>  data <= "11111111";  -- AEA = FF
      when "0101011101011" =>  data <= "11111111";  -- AEB = FF
      when "0101011101100" =>  data <= "11111111";  -- AEC = FF
      when "0101011101101" =>  data <= "11111111";  -- AED = FF
      when "0101011101110" =>  data <= "11111111";  -- AEE = FF
      when "0101011101111" =>  data <= "11111111";  -- AEF = FF
      when "0101011110000" =>  data <= "11111111";  -- AF0 = FF
      when "0101011110001" =>  data <= "11111111";  -- AF1 = FF
      when "0101011110010" =>  data <= "11111111";  -- AF2 = FF
      when "0101011110011" =>  data <= "11111111";  -- AF3 = FF
      when "0101011110100" =>  data <= "11111111";  -- AF4 = FF
      when "0101011110101" =>  data <= "11111111";  -- AF5 = FF
      when "0101011110110" =>  data <= "11111111";  -- AF6 = FF
      when "0101011110111" =>  data <= "11111111";  -- AF7 = FF
      when "0101011111000" =>  data <= "11111111";  -- AF8 = FF
      when "0101011111001" =>  data <= "11111111";  -- AF9 = FF
      when "0101011111010" =>  data <= "11111111";  -- AFA = FF
      when "0101011111011" =>  data <= "11111111";  -- AFB = FF
      when "0101011111100" =>  data <= "11111111";  -- AFC = FF
      when "0101011111101" =>  data <= "11111111";  -- AFD = FF
      when "0101011111110" =>  data <= "11111111";  -- AFE = FF
      when "0101011111111" =>  data <= "11111111";  -- AFF = FF
      when "0101100000000" =>  data <= "11111111";  -- B00 = FF
      when "0101100000001" =>  data <= "11111111";  -- B01 = FF
      when "0101100000010" =>  data <= "11111111";  -- B02 = FF
      when "0101100000011" =>  data <= "11111111";  -- B03 = FF
      when "0101100000100" =>  data <= "11111111";  -- B04 = FF
      when "0101100000101" =>  data <= "11111111";  -- B05 = FF
      when "0101100000110" =>  data <= "11111111";  -- B06 = FF
      when "0101100000111" =>  data <= "11111111";  -- B07 = FF
      when "0101100001000" =>  data <= "11111111";  -- B08 = FF
      when "0101100001001" =>  data <= "11111111";  -- B09 = FF
      when "0101100001010" =>  data <= "11111111";  -- B0A = FF
      when "0101100001011" =>  data <= "11111111";  -- B0B = FF
      when "0101100001100" =>  data <= "11111111";  -- B0C = FF
      when "0101100001101" =>  data <= "11111111";  -- B0D = FF
      when "0101100001110" =>  data <= "11111111";  -- B0E = FF
      when "0101100001111" =>  data <= "11111111";  -- B0F = FF
      when "0101100010000" =>  data <= "11111111";  -- B10 = FF
      when "0101100010001" =>  data <= "11111111";  -- B11 = FF
      when "0101100010010" =>  data <= "11111111";  -- B12 = FF
      when "0101100010011" =>  data <= "11111111";  -- B13 = FF
      when "0101100010100" =>  data <= "11111111";  -- B14 = FF
      when "0101100010101" =>  data <= "11111111";  -- B15 = FF
      when "0101100010110" =>  data <= "11111111";  -- B16 = FF
      when "0101100010111" =>  data <= "11111111";  -- B17 = FF
      when "0101100011000" =>  data <= "11111111";  -- B18 = FF
      when "0101100011001" =>  data <= "11111111";  -- B19 = FF
      when "0101100011010" =>  data <= "11111111";  -- B1A = FF
      when "0101100011011" =>  data <= "11111111";  -- B1B = FF
      when "0101100011100" =>  data <= "11111111";  -- B1C = FF
      when "0101100011101" =>  data <= "11111111";  -- B1D = FF
      when "0101100011110" =>  data <= "11111111";  -- B1E = FF
      when "0101100011111" =>  data <= "11111111";  -- B1F = FF
      when "0101100100000" =>  data <= "11111111";  -- B20 = FF
      when "0101100100001" =>  data <= "11111111";  -- B21 = FF
      when "0101100100010" =>  data <= "11111111";  -- B22 = FF
      when "0101100100011" =>  data <= "11111111";  -- B23 = FF
      when "0101100100100" =>  data <= "11111111";  -- B24 = FF
      when "0101100100101" =>  data <= "11111111";  -- B25 = FF
      when "0101100100110" =>  data <= "11111111";  -- B26 = FF
      when "0101100100111" =>  data <= "11111111";  -- B27 = FF
      when "0101100101000" =>  data <= "11111111";  -- B28 = FF
      when "0101100101001" =>  data <= "11111111";  -- B29 = FF
      when "0101100101010" =>  data <= "11111111";  -- B2A = FF
      when "0101100101011" =>  data <= "11111111";  -- B2B = FF
      when "0101100101100" =>  data <= "11111111";  -- B2C = FF
      when "0101100101101" =>  data <= "11111111";  -- B2D = FF
      when "0101100101110" =>  data <= "11111111";  -- B2E = FF
      when "0101100101111" =>  data <= "11111111";  -- B2F = FF
      when "0101100110000" =>  data <= "11111111";  -- B30 = FF
      when "0101100110001" =>  data <= "11111111";  -- B31 = FF
      when "0101100110010" =>  data <= "11111111";  -- B32 = FF
      when "0101100110011" =>  data <= "11111111";  -- B33 = FF
      when "0101100110100" =>  data <= "11111111";  -- B34 = FF
      when "0101100110101" =>  data <= "11111111";  -- B35 = FF
      when "0101100110110" =>  data <= "11111111";  -- B36 = FF
      when "0101100110111" =>  data <= "11111111";  -- B37 = FF
      when "0101100111000" =>  data <= "11111111";  -- B38 = FF
      when "0101100111001" =>  data <= "11111111";  -- B39 = FF
      when "0101100111010" =>  data <= "11111111";  -- B3A = FF
      when "0101100111011" =>  data <= "11111111";  -- B3B = FF
      when "0101100111100" =>  data <= "11111111";  -- B3C = FF
      when "0101100111101" =>  data <= "11111111";  -- B3D = FF
      when "0101100111110" =>  data <= "11111111";  -- B3E = FF
      when "0101100111111" =>  data <= "11111111";  -- B3F = FF
      when "0101101000000" =>  data <= "11111111";  -- B40 = FF
      when "0101101000001" =>  data <= "11111111";  -- B41 = FF
      when "0101101000010" =>  data <= "11111111";  -- B42 = FF
      when "0101101000011" =>  data <= "11111111";  -- B43 = FF
      when "0101101000100" =>  data <= "11111111";  -- B44 = FF
      when "0101101000101" =>  data <= "11111111";  -- B45 = FF
      when "0101101000110" =>  data <= "11111111";  -- B46 = FF
      when "0101101000111" =>  data <= "11111111";  -- B47 = FF
      when "0101101001000" =>  data <= "11111111";  -- B48 = FF
      when "0101101001001" =>  data <= "11111111";  -- B49 = FF
      when "0101101001010" =>  data <= "11111111";  -- B4A = FF
      when "0101101001011" =>  data <= "11111111";  -- B4B = FF
      when "0101101001100" =>  data <= "11111111";  -- B4C = FF
      when "0101101001101" =>  data <= "11111111";  -- B4D = FF
      when "0101101001110" =>  data <= "11111111";  -- B4E = FF
      when "0101101001111" =>  data <= "11111111";  -- B4F = FF
      when "0101101010000" =>  data <= "11111111";  -- B50 = FF
      when "0101101010001" =>  data <= "11111111";  -- B51 = FF
      when "0101101010010" =>  data <= "11111111";  -- B52 = FF
      when "0101101010011" =>  data <= "11111111";  -- B53 = FF
      when "0101101010100" =>  data <= "11111111";  -- B54 = FF
      when "0101101010101" =>  data <= "11111111";  -- B55 = FF
      when "0101101010110" =>  data <= "11111111";  -- B56 = FF
      when "0101101010111" =>  data <= "11111111";  -- B57 = FF
      when "0101101011000" =>  data <= "11111111";  -- B58 = FF
      when "0101101011001" =>  data <= "11111111";  -- B59 = FF
      when "0101101011010" =>  data <= "11111111";  -- B5A = FF
      when "0101101011011" =>  data <= "11111111";  -- B5B = FF
      when "0101101011100" =>  data <= "11111111";  -- B5C = FF
      when "0101101011101" =>  data <= "11111111";  -- B5D = FF
      when "0101101011110" =>  data <= "11111111";  -- B5E = FF
      when "0101101011111" =>  data <= "11111111";  -- B5F = FF
      when "0101101100000" =>  data <= "11111111";  -- B60 = FF
      when "0101101100001" =>  data <= "11111111";  -- B61 = FF
      when "0101101100010" =>  data <= "11111111";  -- B62 = FF
      when "0101101100011" =>  data <= "11111111";  -- B63 = FF
      when "0101101100100" =>  data <= "11111111";  -- B64 = FF
      when "0101101100101" =>  data <= "11111111";  -- B65 = FF
      when "0101101100110" =>  data <= "11111111";  -- B66 = FF
      when "0101101100111" =>  data <= "11111111";  -- B67 = FF
      when "0101101101000" =>  data <= "11111111";  -- B68 = FF
      when "0101101101001" =>  data <= "11111111";  -- B69 = FF
      when "0101101101010" =>  data <= "11111111";  -- B6A = FF
      when "0101101101011" =>  data <= "11111111";  -- B6B = FF
      when "0101101101100" =>  data <= "11111111";  -- B6C = FF
      when "0101101101101" =>  data <= "11111111";  -- B6D = FF
      when "0101101101110" =>  data <= "11111111";  -- B6E = FF
      when "0101101101111" =>  data <= "11111111";  -- B6F = FF
      when "0101101110000" =>  data <= "11111111";  -- B70 = FF
      when "0101101110001" =>  data <= "11111111";  -- B71 = FF
      when "0101101110010" =>  data <= "11111111";  -- B72 = FF
      when "0101101110011" =>  data <= "11111111";  -- B73 = FF
      when "0101101110100" =>  data <= "11111111";  -- B74 = FF
      when "0101101110101" =>  data <= "11111111";  -- B75 = FF
      when "0101101110110" =>  data <= "11111111";  -- B76 = FF
      when "0101101110111" =>  data <= "11111111";  -- B77 = FF
      when "0101101111000" =>  data <= "11111111";  -- B78 = FF
      when "0101101111001" =>  data <= "11111111";  -- B79 = FF
      when "0101101111010" =>  data <= "11111111";  -- B7A = FF
      when "0101101111011" =>  data <= "11111111";  -- B7B = FF
      when "0101101111100" =>  data <= "11111111";  -- B7C = FF
      when "0101101111101" =>  data <= "11111111";  -- B7D = FF
      when "0101101111110" =>  data <= "11111111";  -- B7E = FF
      when "0101101111111" =>  data <= "11111111";  -- B7F = FF
      when "0101110000000" =>  data <= "11111111";  -- B80 = FF
      when "0101110000001" =>  data <= "11111111";  -- B81 = FF
      when "0101110000010" =>  data <= "11111111";  -- B82 = FF
      when "0101110000011" =>  data <= "11111111";  -- B83 = FF
      when "0101110000100" =>  data <= "11111111";  -- B84 = FF
      when "0101110000101" =>  data <= "11111111";  -- B85 = FF
      when "0101110000110" =>  data <= "11111111";  -- B86 = FF
      when "0101110000111" =>  data <= "11111111";  -- B87 = FF
      when "0101110001000" =>  data <= "11111111";  -- B88 = FF
      when "0101110001001" =>  data <= "11111111";  -- B89 = FF
      when "0101110001010" =>  data <= "11111111";  -- B8A = FF
      when "0101110001011" =>  data <= "11111111";  -- B8B = FF
      when "0101110001100" =>  data <= "11111111";  -- B8C = FF
      when "0101110001101" =>  data <= "11111111";  -- B8D = FF
      when "0101110001110" =>  data <= "11111111";  -- B8E = FF
      when "0101110001111" =>  data <= "11111111";  -- B8F = FF
      when "0101110010000" =>  data <= "11111111";  -- B90 = FF
      when "0101110010001" =>  data <= "11111111";  -- B91 = FF
      when "0101110010010" =>  data <= "11111111";  -- B92 = FF
      when "0101110010011" =>  data <= "11111111";  -- B93 = FF
      when "0101110010100" =>  data <= "11111111";  -- B94 = FF
      when "0101110010101" =>  data <= "11111111";  -- B95 = FF
      when "0101110010110" =>  data <= "11111111";  -- B96 = FF
      when "0101110010111" =>  data <= "11111111";  -- B97 = FF
      when "0101110011000" =>  data <= "11111111";  -- B98 = FF
      when "0101110011001" =>  data <= "11111111";  -- B99 = FF
      when "0101110011010" =>  data <= "11111111";  -- B9A = FF
      when "0101110011011" =>  data <= "11111111";  -- B9B = FF
      when "0101110011100" =>  data <= "11111111";  -- B9C = FF
      when "0101110011101" =>  data <= "11111111";  -- B9D = FF
      when "0101110011110" =>  data <= "11111111";  -- B9E = FF
      when "0101110011111" =>  data <= "11111111";  -- B9F = FF
      when "0101110100000" =>  data <= "11111111";  -- BA0 = FF
      when "0101110100001" =>  data <= "11111111";  -- BA1 = FF
      when "0101110100010" =>  data <= "11111111";  -- BA2 = FF
      when "0101110100011" =>  data <= "11111111";  -- BA3 = FF
      when "0101110100100" =>  data <= "11111111";  -- BA4 = FF
      when "0101110100101" =>  data <= "11111111";  -- BA5 = FF
      when "0101110100110" =>  data <= "11111111";  -- BA6 = FF
      when "0101110100111" =>  data <= "11111111";  -- BA7 = FF
      when "0101110101000" =>  data <= "11111111";  -- BA8 = FF
      when "0101110101001" =>  data <= "11111111";  -- BA9 = FF
      when "0101110101010" =>  data <= "11111111";  -- BAA = FF
      when "0101110101011" =>  data <= "11111111";  -- BAB = FF
      when "0101110101100" =>  data <= "11111111";  -- BAC = FF
      when "0101110101101" =>  data <= "11111111";  -- BAD = FF
      when "0101110101110" =>  data <= "11111111";  -- BAE = FF
      when "0101110101111" =>  data <= "11111111";  -- BAF = FF
      when "0101110110000" =>  data <= "11111111";  -- BB0 = FF
      when "0101110110001" =>  data <= "11111111";  -- BB1 = FF
      when "0101110110010" =>  data <= "11111111";  -- BB2 = FF
      when "0101110110011" =>  data <= "11111111";  -- BB3 = FF
      when "0101110110100" =>  data <= "11111111";  -- BB4 = FF
      when "0101110110101" =>  data <= "11111111";  -- BB5 = FF
      when "0101110110110" =>  data <= "11111111";  -- BB6 = FF
      when "0101110110111" =>  data <= "11111111";  -- BB7 = FF
      when "0101110111000" =>  data <= "11111111";  -- BB8 = FF
      when "0101110111001" =>  data <= "11111111";  -- BB9 = FF
      when "0101110111010" =>  data <= "11111111";  -- BBA = FF
      when "0101110111011" =>  data <= "11111111";  -- BBB = FF
      when "0101110111100" =>  data <= "11111111";  -- BBC = FF
      when "0101110111101" =>  data <= "11111111";  -- BBD = FF
      when "0101110111110" =>  data <= "11111111";  -- BBE = FF
      when "0101110111111" =>  data <= "11111111";  -- BBF = FF
      when "0101111000000" =>  data <= "11111111";  -- BC0 = FF
      when "0101111000001" =>  data <= "11111111";  -- BC1 = FF
      when "0101111000010" =>  data <= "11111111";  -- BC2 = FF
      when "0101111000011" =>  data <= "11111111";  -- BC3 = FF
      when "0101111000100" =>  data <= "11111111";  -- BC4 = FF
      when "0101111000101" =>  data <= "11111111";  -- BC5 = FF
      when "0101111000110" =>  data <= "11111111";  -- BC6 = FF
      when "0101111000111" =>  data <= "11111111";  -- BC7 = FF
      when "0101111001000" =>  data <= "11111111";  -- BC8 = FF
      when "0101111001001" =>  data <= "11111111";  -- BC9 = FF
      when "0101111001010" =>  data <= "11111111";  -- BCA = FF
      when "0101111001011" =>  data <= "11111111";  -- BCB = FF
      when "0101111001100" =>  data <= "11111111";  -- BCC = FF
      when "0101111001101" =>  data <= "11111111";  -- BCD = FF
      when "0101111001110" =>  data <= "11111111";  -- BCE = FF
      when "0101111001111" =>  data <= "11111111";  -- BCF = FF
      when "0101111010000" =>  data <= "11111111";  -- BD0 = FF
      when "0101111010001" =>  data <= "11111111";  -- BD1 = FF
      when "0101111010010" =>  data <= "11111111";  -- BD2 = FF
      when "0101111010011" =>  data <= "11111111";  -- BD3 = FF
      when "0101111010100" =>  data <= "11111111";  -- BD4 = FF
      when "0101111010101" =>  data <= "11111111";  -- BD5 = FF
      when "0101111010110" =>  data <= "11111111";  -- BD6 = FF
      when "0101111010111" =>  data <= "11111111";  -- BD7 = FF
      when "0101111011000" =>  data <= "11111111";  -- BD8 = FF
      when "0101111011001" =>  data <= "11111111";  -- BD9 = FF
      when "0101111011010" =>  data <= "11111111";  -- BDA = FF
      when "0101111011011" =>  data <= "11111111";  -- BDB = FF
      when "0101111011100" =>  data <= "11111111";  -- BDC = FF
      when "0101111011101" =>  data <= "11111111";  -- BDD = FF
      when "0101111011110" =>  data <= "11111111";  -- BDE = FF
      when "0101111011111" =>  data <= "11111111";  -- BDF = FF
      when "0101111100000" =>  data <= "11111111";  -- BE0 = FF
      when "0101111100001" =>  data <= "11111111";  -- BE1 = FF
      when "0101111100010" =>  data <= "11111111";  -- BE2 = FF
      when "0101111100011" =>  data <= "11111111";  -- BE3 = FF
      when "0101111100100" =>  data <= "11111111";  -- BE4 = FF
      when "0101111100101" =>  data <= "11111111";  -- BE5 = FF
      when "0101111100110" =>  data <= "11111111";  -- BE6 = FF
      when "0101111100111" =>  data <= "11111111";  -- BE7 = FF
      when "0101111101000" =>  data <= "11111111";  -- BE8 = FF
      when "0101111101001" =>  data <= "11111111";  -- BE9 = FF
      when "0101111101010" =>  data <= "11111111";  -- BEA = FF
      when "0101111101011" =>  data <= "11111111";  -- BEB = FF
      when "0101111101100" =>  data <= "11111111";  -- BEC = FF
      when "0101111101101" =>  data <= "11111111";  -- BED = FF
      when "0101111101110" =>  data <= "11111111";  -- BEE = FF
      when "0101111101111" =>  data <= "11111111";  -- BEF = FF
      when "0101111110000" =>  data <= "11111111";  -- BF0 = FF
      when "0101111110001" =>  data <= "11111111";  -- BF1 = FF
      when "0101111110010" =>  data <= "11111111";  -- BF2 = FF
      when "0101111110011" =>  data <= "11111111";  -- BF3 = FF
      when "0101111110100" =>  data <= "11111111";  -- BF4 = FF
      when "0101111110101" =>  data <= "11111111";  -- BF5 = FF
      when "0101111110110" =>  data <= "11111111";  -- BF6 = FF
      when "0101111110111" =>  data <= "11111111";  -- BF7 = FF
      when "0101111111000" =>  data <= "11111111";  -- BF8 = FF
      when "0101111111001" =>  data <= "11111111";  -- BF9 = FF
      when "0101111111010" =>  data <= "11111111";  -- BFA = FF
      when "0101111111011" =>  data <= "11111111";  -- BFB = FF
      when "0101111111100" =>  data <= "11111111";  -- BFC = FF
      when "0101111111101" =>  data <= "11111111";  -- BFD = FF
      when "0101111111110" =>  data <= "11111111";  -- BFE = FF
      when "0101111111111" =>  data <= "11111111";  -- BFF = FF
      when "0110000000000" =>  data <= "11111111";  -- C00 = FF
      when "0110000000001" =>  data <= "11111111";  -- C01 = FF
      when "0110000000010" =>  data <= "11111111";  -- C02 = FF
      when "0110000000011" =>  data <= "11111111";  -- C03 = FF
      when "0110000000100" =>  data <= "11111111";  -- C04 = FF
      when "0110000000101" =>  data <= "11111111";  -- C05 = FF
      when "0110000000110" =>  data <= "11111111";  -- C06 = FF
      when "0110000000111" =>  data <= "11111111";  -- C07 = FF
      when "0110000001000" =>  data <= "11111111";  -- C08 = FF
      when "0110000001001" =>  data <= "11111111";  -- C09 = FF
      when "0110000001010" =>  data <= "11111111";  -- C0A = FF
      when "0110000001011" =>  data <= "11111111";  -- C0B = FF
      when "0110000001100" =>  data <= "11111111";  -- C0C = FF
      when "0110000001101" =>  data <= "11111111";  -- C0D = FF
      when "0110000001110" =>  data <= "11111111";  -- C0E = FF
      when "0110000001111" =>  data <= "11111111";  -- C0F = FF
      when "0110000010000" =>  data <= "11111111";  -- C10 = FF
      when "0110000010001" =>  data <= "11111111";  -- C11 = FF
      when "0110000010010" =>  data <= "11111111";  -- C12 = FF
      when "0110000010011" =>  data <= "11111111";  -- C13 = FF
      when "0110000010100" =>  data <= "11111111";  -- C14 = FF
      when "0110000010101" =>  data <= "11111111";  -- C15 = FF
      when "0110000010110" =>  data <= "11111111";  -- C16 = FF
      when "0110000010111" =>  data <= "11111111";  -- C17 = FF
      when "0110000011000" =>  data <= "11111111";  -- C18 = FF
      when "0110000011001" =>  data <= "11111111";  -- C19 = FF
      when "0110000011010" =>  data <= "11111111";  -- C1A = FF
      when "0110000011011" =>  data <= "11111111";  -- C1B = FF
      when "0110000011100" =>  data <= "11111111";  -- C1C = FF
      when "0110000011101" =>  data <= "11111111";  -- C1D = FF
      when "0110000011110" =>  data <= "11111111";  -- C1E = FF
      when "0110000011111" =>  data <= "11111111";  -- C1F = FF
      when "0110000100000" =>  data <= "11111111";  -- C20 = FF
      when "0110000100001" =>  data <= "11111111";  -- C21 = FF
      when "0110000100010" =>  data <= "11111111";  -- C22 = FF
      when "0110000100011" =>  data <= "11111111";  -- C23 = FF
      when "0110000100100" =>  data <= "11111111";  -- C24 = FF
      when "0110000100101" =>  data <= "11111111";  -- C25 = FF
      when "0110000100110" =>  data <= "11111111";  -- C26 = FF
      when "0110000100111" =>  data <= "11111111";  -- C27 = FF
      when "0110000101000" =>  data <= "11111111";  -- C28 = FF
      when "0110000101001" =>  data <= "11111111";  -- C29 = FF
      when "0110000101010" =>  data <= "11111111";  -- C2A = FF
      when "0110000101011" =>  data <= "11111111";  -- C2B = FF
      when "0110000101100" =>  data <= "11111111";  -- C2C = FF
      when "0110000101101" =>  data <= "11111111";  -- C2D = FF
      when "0110000101110" =>  data <= "11111111";  -- C2E = FF
      when "0110000101111" =>  data <= "11111111";  -- C2F = FF
      when "0110000110000" =>  data <= "11111111";  -- C30 = FF
      when "0110000110001" =>  data <= "11111111";  -- C31 = FF
      when "0110000110010" =>  data <= "11111111";  -- C32 = FF
      when "0110000110011" =>  data <= "11111111";  -- C33 = FF
      when "0110000110100" =>  data <= "11111111";  -- C34 = FF
      when "0110000110101" =>  data <= "11111111";  -- C35 = FF
      when "0110000110110" =>  data <= "11111111";  -- C36 = FF
      when "0110000110111" =>  data <= "11111111";  -- C37 = FF
      when "0110000111000" =>  data <= "11111111";  -- C38 = FF
      when "0110000111001" =>  data <= "11111111";  -- C39 = FF
      when "0110000111010" =>  data <= "11111111";  -- C3A = FF
      when "0110000111011" =>  data <= "11111111";  -- C3B = FF
      when "0110000111100" =>  data <= "11111111";  -- C3C = FF
      when "0110000111101" =>  data <= "11111111";  -- C3D = FF
      when "0110000111110" =>  data <= "11111111";  -- C3E = FF
      when "0110000111111" =>  data <= "11111111";  -- C3F = FF
      when "0110001000000" =>  data <= "11111111";  -- C40 = FF
      when "0110001000001" =>  data <= "11111111";  -- C41 = FF
      when "0110001000010" =>  data <= "11111111";  -- C42 = FF
      when "0110001000011" =>  data <= "11111111";  -- C43 = FF
      when "0110001000100" =>  data <= "11111111";  -- C44 = FF
      when "0110001000101" =>  data <= "11111111";  -- C45 = FF
      when "0110001000110" =>  data <= "11111111";  -- C46 = FF
      when "0110001000111" =>  data <= "11111111";  -- C47 = FF
      when "0110001001000" =>  data <= "11111111";  -- C48 = FF
      when "0110001001001" =>  data <= "11111111";  -- C49 = FF
      when "0110001001010" =>  data <= "11111111";  -- C4A = FF
      when "0110001001011" =>  data <= "11111111";  -- C4B = FF
      when "0110001001100" =>  data <= "11111111";  -- C4C = FF
      when "0110001001101" =>  data <= "11111111";  -- C4D = FF
      when "0110001001110" =>  data <= "11111111";  -- C4E = FF
      when "0110001001111" =>  data <= "11111111";  -- C4F = FF
      when "0110001010000" =>  data <= "11111111";  -- C50 = FF
      when "0110001010001" =>  data <= "11111111";  -- C51 = FF
      when "0110001010010" =>  data <= "11111111";  -- C52 = FF
      when "0110001010011" =>  data <= "11111111";  -- C53 = FF
      when "0110001010100" =>  data <= "11111111";  -- C54 = FF
      when "0110001010101" =>  data <= "11111111";  -- C55 = FF
      when "0110001010110" =>  data <= "11111111";  -- C56 = FF
      when "0110001010111" =>  data <= "11111111";  -- C57 = FF
      when "0110001011000" =>  data <= "11111111";  -- C58 = FF
      when "0110001011001" =>  data <= "11111111";  -- C59 = FF
      when "0110001011010" =>  data <= "11111111";  -- C5A = FF
      when "0110001011011" =>  data <= "11111111";  -- C5B = FF
      when "0110001011100" =>  data <= "11111111";  -- C5C = FF
      when "0110001011101" =>  data <= "11111111";  -- C5D = FF
      when "0110001011110" =>  data <= "11111111";  -- C5E = FF
      when "0110001011111" =>  data <= "11111111";  -- C5F = FF
      when "0110001100000" =>  data <= "11111111";  -- C60 = FF
      when "0110001100001" =>  data <= "11111111";  -- C61 = FF
      when "0110001100010" =>  data <= "11111111";  -- C62 = FF
      when "0110001100011" =>  data <= "11111111";  -- C63 = FF
      when "0110001100100" =>  data <= "11111111";  -- C64 = FF
      when "0110001100101" =>  data <= "11111111";  -- C65 = FF
      when "0110001100110" =>  data <= "11111111";  -- C66 = FF
      when "0110001100111" =>  data <= "11111111";  -- C67 = FF
      when "0110001101000" =>  data <= "11111111";  -- C68 = FF
      when "0110001101001" =>  data <= "11111111";  -- C69 = FF
      when "0110001101010" =>  data <= "11111111";  -- C6A = FF
      when "0110001101011" =>  data <= "11111111";  -- C6B = FF
      when "0110001101100" =>  data <= "11111111";  -- C6C = FF
      when "0110001101101" =>  data <= "11111111";  -- C6D = FF
      when "0110001101110" =>  data <= "11111111";  -- C6E = FF
      when "0110001101111" =>  data <= "11111111";  -- C6F = FF
      when "0110001110000" =>  data <= "11111111";  -- C70 = FF
      when "0110001110001" =>  data <= "11111111";  -- C71 = FF
      when "0110001110010" =>  data <= "11111111";  -- C72 = FF
      when "0110001110011" =>  data <= "11111111";  -- C73 = FF
      when "0110001110100" =>  data <= "11111111";  -- C74 = FF
      when "0110001110101" =>  data <= "11111111";  -- C75 = FF
      when "0110001110110" =>  data <= "11111111";  -- C76 = FF
      when "0110001110111" =>  data <= "11111111";  -- C77 = FF
      when "0110001111000" =>  data <= "11111111";  -- C78 = FF
      when "0110001111001" =>  data <= "11111111";  -- C79 = FF
      when "0110001111010" =>  data <= "11111111";  -- C7A = FF
      when "0110001111011" =>  data <= "11111111";  -- C7B = FF
      when "0110001111100" =>  data <= "11111111";  -- C7C = FF
      when "0110001111101" =>  data <= "11111111";  -- C7D = FF
      when "0110001111110" =>  data <= "11111111";  -- C7E = FF
      when "0110001111111" =>  data <= "11111111";  -- C7F = FF
      when "0110010000000" =>  data <= "11111111";  -- C80 = FF
      when "0110010000001" =>  data <= "11111111";  -- C81 = FF
      when "0110010000010" =>  data <= "11111111";  -- C82 = FF
      when "0110010000011" =>  data <= "11111111";  -- C83 = FF
      when "0110010000100" =>  data <= "11111111";  -- C84 = FF
      when "0110010000101" =>  data <= "11111111";  -- C85 = FF
      when "0110010000110" =>  data <= "11111111";  -- C86 = FF
      when "0110010000111" =>  data <= "11111111";  -- C87 = FF
      when "0110010001000" =>  data <= "11111111";  -- C88 = FF
      when "0110010001001" =>  data <= "11111111";  -- C89 = FF
      when "0110010001010" =>  data <= "11111111";  -- C8A = FF
      when "0110010001011" =>  data <= "11111111";  -- C8B = FF
      when "0110010001100" =>  data <= "11111111";  -- C8C = FF
      when "0110010001101" =>  data <= "11111111";  -- C8D = FF
      when "0110010001110" =>  data <= "11111111";  -- C8E = FF
      when "0110010001111" =>  data <= "11111111";  -- C8F = FF
      when "0110010010000" =>  data <= "11111111";  -- C90 = FF
      when "0110010010001" =>  data <= "11111111";  -- C91 = FF
      when "0110010010010" =>  data <= "11111111";  -- C92 = FF
      when "0110010010011" =>  data <= "11111111";  -- C93 = FF
      when "0110010010100" =>  data <= "11111111";  -- C94 = FF
      when "0110010010101" =>  data <= "11111111";  -- C95 = FF
      when "0110010010110" =>  data <= "11111111";  -- C96 = FF
      when "0110010010111" =>  data <= "11111111";  -- C97 = FF
      when "0110010011000" =>  data <= "11111111";  -- C98 = FF
      when "0110010011001" =>  data <= "11111111";  -- C99 = FF
      when "0110010011010" =>  data <= "11111111";  -- C9A = FF
      when "0110010011011" =>  data <= "11111111";  -- C9B = FF
      when "0110010011100" =>  data <= "11111111";  -- C9C = FF
      when "0110010011101" =>  data <= "11111111";  -- C9D = FF
      when "0110010011110" =>  data <= "11111111";  -- C9E = FF
      when "0110010011111" =>  data <= "11111111";  -- C9F = FF
      when "0110010100000" =>  data <= "11111111";  -- CA0 = FF
      when "0110010100001" =>  data <= "11111111";  -- CA1 = FF
      when "0110010100010" =>  data <= "11111111";  -- CA2 = FF
      when "0110010100011" =>  data <= "11111111";  -- CA3 = FF
      when "0110010100100" =>  data <= "11111111";  -- CA4 = FF
      when "0110010100101" =>  data <= "11111111";  -- CA5 = FF
      when "0110010100110" =>  data <= "11111111";  -- CA6 = FF
      when "0110010100111" =>  data <= "11111111";  -- CA7 = FF
      when "0110010101000" =>  data <= "11111111";  -- CA8 = FF
      when "0110010101001" =>  data <= "11111111";  -- CA9 = FF
      when "0110010101010" =>  data <= "11111111";  -- CAA = FF
      when "0110010101011" =>  data <= "11111111";  -- CAB = FF
      when "0110010101100" =>  data <= "11111111";  -- CAC = FF
      when "0110010101101" =>  data <= "11111111";  -- CAD = FF
      when "0110010101110" =>  data <= "11111111";  -- CAE = FF
      when "0110010101111" =>  data <= "11111111";  -- CAF = FF
      when "0110010110000" =>  data <= "11111111";  -- CB0 = FF
      when "0110010110001" =>  data <= "11111111";  -- CB1 = FF
      when "0110010110010" =>  data <= "11111111";  -- CB2 = FF
      when "0110010110011" =>  data <= "11111111";  -- CB3 = FF
      when "0110010110100" =>  data <= "11111111";  -- CB4 = FF
      when "0110010110101" =>  data <= "11111111";  -- CB5 = FF
      when "0110010110110" =>  data <= "11111111";  -- CB6 = FF
      when "0110010110111" =>  data <= "11111111";  -- CB7 = FF
      when "0110010111000" =>  data <= "11111111";  -- CB8 = FF
      when "0110010111001" =>  data <= "11111111";  -- CB9 = FF
      when "0110010111010" =>  data <= "11111111";  -- CBA = FF
      when "0110010111011" =>  data <= "11111111";  -- CBB = FF
      when "0110010111100" =>  data <= "11111111";  -- CBC = FF
      when "0110010111101" =>  data <= "11111111";  -- CBD = FF
      when "0110010111110" =>  data <= "11111111";  -- CBE = FF
      when "0110010111111" =>  data <= "11111111";  -- CBF = FF
      when "0110011000000" =>  data <= "11111111";  -- CC0 = FF
      when "0110011000001" =>  data <= "11111111";  -- CC1 = FF
      when "0110011000010" =>  data <= "11111111";  -- CC2 = FF
      when "0110011000011" =>  data <= "11111111";  -- CC3 = FF
      when "0110011000100" =>  data <= "11111111";  -- CC4 = FF
      when "0110011000101" =>  data <= "11111111";  -- CC5 = FF
      when "0110011000110" =>  data <= "11111111";  -- CC6 = FF
      when "0110011000111" =>  data <= "11111111";  -- CC7 = FF
      when "0110011001000" =>  data <= "11111111";  -- CC8 = FF
      when "0110011001001" =>  data <= "11111111";  -- CC9 = FF
      when "0110011001010" =>  data <= "11111111";  -- CCA = FF
      when "0110011001011" =>  data <= "11111111";  -- CCB = FF
      when "0110011001100" =>  data <= "11111111";  -- CCC = FF
      when "0110011001101" =>  data <= "11111111";  -- CCD = FF
      when "0110011001110" =>  data <= "11111111";  -- CCE = FF
      when "0110011001111" =>  data <= "11111111";  -- CCF = FF
      when "0110011010000" =>  data <= "11111111";  -- CD0 = FF
      when "0110011010001" =>  data <= "11111111";  -- CD1 = FF
      when "0110011010010" =>  data <= "11111111";  -- CD2 = FF
      when "0110011010011" =>  data <= "11111111";  -- CD3 = FF
      when "0110011010100" =>  data <= "11111111";  -- CD4 = FF
      when "0110011010101" =>  data <= "11111111";  -- CD5 = FF
      when "0110011010110" =>  data <= "11111111";  -- CD6 = FF
      when "0110011010111" =>  data <= "11111111";  -- CD7 = FF
      when "0110011011000" =>  data <= "11111111";  -- CD8 = FF
      when "0110011011001" =>  data <= "11111111";  -- CD9 = FF
      when "0110011011010" =>  data <= "11111111";  -- CDA = FF
      when "0110011011011" =>  data <= "11111111";  -- CDB = FF
      when "0110011011100" =>  data <= "11111111";  -- CDC = FF
      when "0110011011101" =>  data <= "11111111";  -- CDD = FF
      when "0110011011110" =>  data <= "11111111";  -- CDE = FF
      when "0110011011111" =>  data <= "11111111";  -- CDF = FF
      when "0110011100000" =>  data <= "11111111";  -- CE0 = FF
      when "0110011100001" =>  data <= "11111111";  -- CE1 = FF
      when "0110011100010" =>  data <= "11111111";  -- CE2 = FF
      when "0110011100011" =>  data <= "11111111";  -- CE3 = FF
      when "0110011100100" =>  data <= "11111111";  -- CE4 = FF
      when "0110011100101" =>  data <= "11111111";  -- CE5 = FF
      when "0110011100110" =>  data <= "11111111";  -- CE6 = FF
      when "0110011100111" =>  data <= "11111111";  -- CE7 = FF
      when "0110011101000" =>  data <= "11111111";  -- CE8 = FF
      when "0110011101001" =>  data <= "11111111";  -- CE9 = FF
      when "0110011101010" =>  data <= "11111111";  -- CEA = FF
      when "0110011101011" =>  data <= "11111111";  -- CEB = FF
      when "0110011101100" =>  data <= "11111111";  -- CEC = FF
      when "0110011101101" =>  data <= "11111111";  -- CED = FF
      when "0110011101110" =>  data <= "11111111";  -- CEE = FF
      when "0110011101111" =>  data <= "11111111";  -- CEF = FF
      when "0110011110000" =>  data <= "11111111";  -- CF0 = FF
      when "0110011110001" =>  data <= "11111111";  -- CF1 = FF
      when "0110011110010" =>  data <= "11111111";  -- CF2 = FF
      when "0110011110011" =>  data <= "11111111";  -- CF3 = FF
      when "0110011110100" =>  data <= "11111111";  -- CF4 = FF
      when "0110011110101" =>  data <= "11111111";  -- CF5 = FF
      when "0110011110110" =>  data <= "11111111";  -- CF6 = FF
      when "0110011110111" =>  data <= "11111111";  -- CF7 = FF
      when "0110011111000" =>  data <= "11111111";  -- CF8 = FF
      when "0110011111001" =>  data <= "11111111";  -- CF9 = FF
      when "0110011111010" =>  data <= "11111111";  -- CFA = FF
      when "0110011111011" =>  data <= "11111111";  -- CFB = FF
      when "0110011111100" =>  data <= "11111111";  -- CFC = FF
      when "0110011111101" =>  data <= "11111111";  -- CFD = FF
      when "0110011111110" =>  data <= "11111111";  -- CFE = FF
      when "0110011111111" =>  data <= "11111111";  -- CFF = FF
      when "0110100000000" =>  data <= "11111111";  -- D00 = FF
      when "0110100000001" =>  data <= "11111111";  -- D01 = FF
      when "0110100000010" =>  data <= "11111111";  -- D02 = FF
      when "0110100000011" =>  data <= "11111111";  -- D03 = FF
      when "0110100000100" =>  data <= "11111111";  -- D04 = FF
      when "0110100000101" =>  data <= "11111111";  -- D05 = FF
      when "0110100000110" =>  data <= "11111111";  -- D06 = FF
      when "0110100000111" =>  data <= "11111111";  -- D07 = FF
      when "0110100001000" =>  data <= "11111111";  -- D08 = FF
      when "0110100001001" =>  data <= "11111111";  -- D09 = FF
      when "0110100001010" =>  data <= "11111111";  -- D0A = FF
      when "0110100001011" =>  data <= "11111111";  -- D0B = FF
      when "0110100001100" =>  data <= "11111111";  -- D0C = FF
      when "0110100001101" =>  data <= "11111111";  -- D0D = FF
      when "0110100001110" =>  data <= "11111111";  -- D0E = FF
      when "0110100001111" =>  data <= "11111111";  -- D0F = FF
      when "0110100010000" =>  data <= "11111111";  -- D10 = FF
      when "0110100010001" =>  data <= "11111111";  -- D11 = FF
      when "0110100010010" =>  data <= "11111111";  -- D12 = FF
      when "0110100010011" =>  data <= "11111111";  -- D13 = FF
      when "0110100010100" =>  data <= "11111111";  -- D14 = FF
      when "0110100010101" =>  data <= "11111111";  -- D15 = FF
      when "0110100010110" =>  data <= "11111111";  -- D16 = FF
      when "0110100010111" =>  data <= "11111111";  -- D17 = FF
      when "0110100011000" =>  data <= "11111111";  -- D18 = FF
      when "0110100011001" =>  data <= "11111111";  -- D19 = FF
      when "0110100011010" =>  data <= "11111111";  -- D1A = FF
      when "0110100011011" =>  data <= "11111111";  -- D1B = FF
      when "0110100011100" =>  data <= "11111111";  -- D1C = FF
      when "0110100011101" =>  data <= "11111111";  -- D1D = FF
      when "0110100011110" =>  data <= "11111111";  -- D1E = FF
      when "0110100011111" =>  data <= "11111111";  -- D1F = FF
      when "0110100100000" =>  data <= "11111111";  -- D20 = FF
      when "0110100100001" =>  data <= "11111111";  -- D21 = FF
      when "0110100100010" =>  data <= "11111111";  -- D22 = FF
      when "0110100100011" =>  data <= "11111111";  -- D23 = FF
      when "0110100100100" =>  data <= "11111111";  -- D24 = FF
      when "0110100100101" =>  data <= "11111111";  -- D25 = FF
      when "0110100100110" =>  data <= "11111111";  -- D26 = FF
      when "0110100100111" =>  data <= "11111111";  -- D27 = FF
      when "0110100101000" =>  data <= "11111111";  -- D28 = FF
      when "0110100101001" =>  data <= "11111111";  -- D29 = FF
      when "0110100101010" =>  data <= "11111111";  -- D2A = FF
      when "0110100101011" =>  data <= "11111111";  -- D2B = FF
      when "0110100101100" =>  data <= "11111111";  -- D2C = FF
      when "0110100101101" =>  data <= "11111111";  -- D2D = FF
      when "0110100101110" =>  data <= "11111111";  -- D2E = FF
      when "0110100101111" =>  data <= "11111111";  -- D2F = FF
      when "0110100110000" =>  data <= "11111111";  -- D30 = FF
      when "0110100110001" =>  data <= "11111111";  -- D31 = FF
      when "0110100110010" =>  data <= "11111111";  -- D32 = FF
      when "0110100110011" =>  data <= "11111111";  -- D33 = FF
      when "0110100110100" =>  data <= "11111111";  -- D34 = FF
      when "0110100110101" =>  data <= "11111111";  -- D35 = FF
      when "0110100110110" =>  data <= "11111111";  -- D36 = FF
      when "0110100110111" =>  data <= "11111111";  -- D37 = FF
      when "0110100111000" =>  data <= "11111111";  -- D38 = FF
      when "0110100111001" =>  data <= "11111111";  -- D39 = FF
      when "0110100111010" =>  data <= "11111111";  -- D3A = FF
      when "0110100111011" =>  data <= "11111111";  -- D3B = FF
      when "0110100111100" =>  data <= "11111111";  -- D3C = FF
      when "0110100111101" =>  data <= "11111111";  -- D3D = FF
      when "0110100111110" =>  data <= "11111111";  -- D3E = FF
      when "0110100111111" =>  data <= "11111111";  -- D3F = FF
      when "0110101000000" =>  data <= "11111111";  -- D40 = FF
      when "0110101000001" =>  data <= "11111111";  -- D41 = FF
      when "0110101000010" =>  data <= "11111111";  -- D42 = FF
      when "0110101000011" =>  data <= "11111111";  -- D43 = FF
      when "0110101000100" =>  data <= "11111111";  -- D44 = FF
      when "0110101000101" =>  data <= "11111111";  -- D45 = FF
      when "0110101000110" =>  data <= "11111111";  -- D46 = FF
      when "0110101000111" =>  data <= "11111111";  -- D47 = FF
      when "0110101001000" =>  data <= "11111111";  -- D48 = FF
      when "0110101001001" =>  data <= "11111111";  -- D49 = FF
      when "0110101001010" =>  data <= "11111111";  -- D4A = FF
      when "0110101001011" =>  data <= "11111111";  -- D4B = FF
      when "0110101001100" =>  data <= "11111111";  -- D4C = FF
      when "0110101001101" =>  data <= "11111111";  -- D4D = FF
      when "0110101001110" =>  data <= "11111111";  -- D4E = FF
      when "0110101001111" =>  data <= "11111111";  -- D4F = FF
      when "0110101010000" =>  data <= "11111111";  -- D50 = FF
      when "0110101010001" =>  data <= "11111111";  -- D51 = FF
      when "0110101010010" =>  data <= "11111111";  -- D52 = FF
      when "0110101010011" =>  data <= "11111111";  -- D53 = FF
      when "0110101010100" =>  data <= "11111111";  -- D54 = FF
      when "0110101010101" =>  data <= "11111111";  -- D55 = FF
      when "0110101010110" =>  data <= "11111111";  -- D56 = FF
      when "0110101010111" =>  data <= "11111111";  -- D57 = FF
      when "0110101011000" =>  data <= "11111111";  -- D58 = FF
      when "0110101011001" =>  data <= "11111111";  -- D59 = FF
      when "0110101011010" =>  data <= "11111111";  -- D5A = FF
      when "0110101011011" =>  data <= "11111111";  -- D5B = FF
      when "0110101011100" =>  data <= "11111111";  -- D5C = FF
      when "0110101011101" =>  data <= "11111111";  -- D5D = FF
      when "0110101011110" =>  data <= "11111111";  -- D5E = FF
      when "0110101011111" =>  data <= "11111111";  -- D5F = FF
      when "0110101100000" =>  data <= "11111111";  -- D60 = FF
      when "0110101100001" =>  data <= "11111111";  -- D61 = FF
      when "0110101100010" =>  data <= "11111111";  -- D62 = FF
      when "0110101100011" =>  data <= "11111111";  -- D63 = FF
      when "0110101100100" =>  data <= "11111111";  -- D64 = FF
      when "0110101100101" =>  data <= "11111111";  -- D65 = FF
      when "0110101100110" =>  data <= "11111111";  -- D66 = FF
      when "0110101100111" =>  data <= "11111111";  -- D67 = FF
      when "0110101101000" =>  data <= "11111111";  -- D68 = FF
      when "0110101101001" =>  data <= "11111111";  -- D69 = FF
      when "0110101101010" =>  data <= "11111111";  -- D6A = FF
      when "0110101101011" =>  data <= "11111111";  -- D6B = FF
      when "0110101101100" =>  data <= "11111111";  -- D6C = FF
      when "0110101101101" =>  data <= "11111111";  -- D6D = FF
      when "0110101101110" =>  data <= "11111111";  -- D6E = FF
      when "0110101101111" =>  data <= "11111111";  -- D6F = FF
      when "0110101110000" =>  data <= "11111111";  -- D70 = FF
      when "0110101110001" =>  data <= "11111111";  -- D71 = FF
      when "0110101110010" =>  data <= "11111111";  -- D72 = FF
      when "0110101110011" =>  data <= "11111111";  -- D73 = FF
      when "0110101110100" =>  data <= "11111111";  -- D74 = FF
      when "0110101110101" =>  data <= "11111111";  -- D75 = FF
      when "0110101110110" =>  data <= "11111111";  -- D76 = FF
      when "0110101110111" =>  data <= "11111111";  -- D77 = FF
      when "0110101111000" =>  data <= "11111111";  -- D78 = FF
      when "0110101111001" =>  data <= "11111111";  -- D79 = FF
      when "0110101111010" =>  data <= "11111111";  -- D7A = FF
      when "0110101111011" =>  data <= "11111111";  -- D7B = FF
      when "0110101111100" =>  data <= "11111111";  -- D7C = FF
      when "0110101111101" =>  data <= "11111111";  -- D7D = FF
      when "0110101111110" =>  data <= "11111111";  -- D7E = FF
      when "0110101111111" =>  data <= "11111111";  -- D7F = FF
      when "0110110000000" =>  data <= "11111111";  -- D80 = FF
      when "0110110000001" =>  data <= "11111111";  -- D81 = FF
      when "0110110000010" =>  data <= "11111111";  -- D82 = FF
      when "0110110000011" =>  data <= "11111111";  -- D83 = FF
      when "0110110000100" =>  data <= "11111111";  -- D84 = FF
      when "0110110000101" =>  data <= "11111111";  -- D85 = FF
      when "0110110000110" =>  data <= "11111111";  -- D86 = FF
      when "0110110000111" =>  data <= "11111111";  -- D87 = FF
      when "0110110001000" =>  data <= "11111111";  -- D88 = FF
      when "0110110001001" =>  data <= "11111111";  -- D89 = FF
      when "0110110001010" =>  data <= "11111111";  -- D8A = FF
      when "0110110001011" =>  data <= "11111111";  -- D8B = FF
      when "0110110001100" =>  data <= "11111111";  -- D8C = FF
      when "0110110001101" =>  data <= "11111111";  -- D8D = FF
      when "0110110001110" =>  data <= "11111111";  -- D8E = FF
      when "0110110001111" =>  data <= "11111111";  -- D8F = FF
      when "0110110010000" =>  data <= "11111111";  -- D90 = FF
      when "0110110010001" =>  data <= "11111111";  -- D91 = FF
      when "0110110010010" =>  data <= "11111111";  -- D92 = FF
      when "0110110010011" =>  data <= "11111111";  -- D93 = FF
      when "0110110010100" =>  data <= "11111111";  -- D94 = FF
      when "0110110010101" =>  data <= "11111111";  -- D95 = FF
      when "0110110010110" =>  data <= "11111111";  -- D96 = FF
      when "0110110010111" =>  data <= "11111111";  -- D97 = FF
      when "0110110011000" =>  data <= "11111111";  -- D98 = FF
      when "0110110011001" =>  data <= "11111111";  -- D99 = FF
      when "0110110011010" =>  data <= "11111111";  -- D9A = FF
      when "0110110011011" =>  data <= "11111111";  -- D9B = FF
      when "0110110011100" =>  data <= "11111111";  -- D9C = FF
      when "0110110011101" =>  data <= "11111111";  -- D9D = FF
      when "0110110011110" =>  data <= "11111111";  -- D9E = FF
      when "0110110011111" =>  data <= "11111111";  -- D9F = FF
      when "0110110100000" =>  data <= "11111111";  -- DA0 = FF
      when "0110110100001" =>  data <= "11111111";  -- DA1 = FF
      when "0110110100010" =>  data <= "11111111";  -- DA2 = FF
      when "0110110100011" =>  data <= "11111111";  -- DA3 = FF
      when "0110110100100" =>  data <= "11111111";  -- DA4 = FF
      when "0110110100101" =>  data <= "11111111";  -- DA5 = FF
      when "0110110100110" =>  data <= "11111111";  -- DA6 = FF
      when "0110110100111" =>  data <= "11111111";  -- DA7 = FF
      when "0110110101000" =>  data <= "11111111";  -- DA8 = FF
      when "0110110101001" =>  data <= "11111111";  -- DA9 = FF
      when "0110110101010" =>  data <= "11111111";  -- DAA = FF
      when "0110110101011" =>  data <= "11111111";  -- DAB = FF
      when "0110110101100" =>  data <= "11111111";  -- DAC = FF
      when "0110110101101" =>  data <= "11111111";  -- DAD = FF
      when "0110110101110" =>  data <= "11111111";  -- DAE = FF
      when "0110110101111" =>  data <= "11111111";  -- DAF = FF
      when "0110110110000" =>  data <= "11111111";  -- DB0 = FF
      when "0110110110001" =>  data <= "11111111";  -- DB1 = FF
      when "0110110110010" =>  data <= "11111111";  -- DB2 = FF
      when "0110110110011" =>  data <= "11111111";  -- DB3 = FF
      when "0110110110100" =>  data <= "11111111";  -- DB4 = FF
      when "0110110110101" =>  data <= "11111111";  -- DB5 = FF
      when "0110110110110" =>  data <= "11111111";  -- DB6 = FF
      when "0110110110111" =>  data <= "11111111";  -- DB7 = FF
      when "0110110111000" =>  data <= "11111111";  -- DB8 = FF
      when "0110110111001" =>  data <= "11111111";  -- DB9 = FF
      when "0110110111010" =>  data <= "11111111";  -- DBA = FF
      when "0110110111011" =>  data <= "11111111";  -- DBB = FF
      when "0110110111100" =>  data <= "11111111";  -- DBC = FF
      when "0110110111101" =>  data <= "11111111";  -- DBD = FF
      when "0110110111110" =>  data <= "11111111";  -- DBE = FF
      when "0110110111111" =>  data <= "11111111";  -- DBF = FF
      when "0110111000000" =>  data <= "11111111";  -- DC0 = FF
      when "0110111000001" =>  data <= "11111111";  -- DC1 = FF
      when "0110111000010" =>  data <= "11111111";  -- DC2 = FF
      when "0110111000011" =>  data <= "11111111";  -- DC3 = FF
      when "0110111000100" =>  data <= "11111111";  -- DC4 = FF
      when "0110111000101" =>  data <= "11111111";  -- DC5 = FF
      when "0110111000110" =>  data <= "11111111";  -- DC6 = FF
      when "0110111000111" =>  data <= "11111111";  -- DC7 = FF
      when "0110111001000" =>  data <= "11111111";  -- DC8 = FF
      when "0110111001001" =>  data <= "11111111";  -- DC9 = FF
      when "0110111001010" =>  data <= "11111111";  -- DCA = FF
      when "0110111001011" =>  data <= "11111111";  -- DCB = FF
      when "0110111001100" =>  data <= "11111111";  -- DCC = FF
      when "0110111001101" =>  data <= "11111111";  -- DCD = FF
      when "0110111001110" =>  data <= "11111111";  -- DCE = FF
      when "0110111001111" =>  data <= "11111111";  -- DCF = FF
      when "0110111010000" =>  data <= "11111111";  -- DD0 = FF
      when "0110111010001" =>  data <= "11111111";  -- DD1 = FF
      when "0110111010010" =>  data <= "11111111";  -- DD2 = FF
      when "0110111010011" =>  data <= "11111111";  -- DD3 = FF
      when "0110111010100" =>  data <= "11111111";  -- DD4 = FF
      when "0110111010101" =>  data <= "11111111";  -- DD5 = FF
      when "0110111010110" =>  data <= "11111111";  -- DD6 = FF
      when "0110111010111" =>  data <= "11111111";  -- DD7 = FF
      when "0110111011000" =>  data <= "11111111";  -- DD8 = FF
      when "0110111011001" =>  data <= "11111111";  -- DD9 = FF
      when "0110111011010" =>  data <= "11111111";  -- DDA = FF
      when "0110111011011" =>  data <= "11111111";  -- DDB = FF
      when "0110111011100" =>  data <= "11111111";  -- DDC = FF
      when "0110111011101" =>  data <= "11111111";  -- DDD = FF
      when "0110111011110" =>  data <= "11111111";  -- DDE = FF
      when "0110111011111" =>  data <= "11111111";  -- DDF = FF
      when "0110111100000" =>  data <= "11111111";  -- DE0 = FF
      when "0110111100001" =>  data <= "11111111";  -- DE1 = FF
      when "0110111100010" =>  data <= "11111111";  -- DE2 = FF
      when "0110111100011" =>  data <= "11111111";  -- DE3 = FF
      when "0110111100100" =>  data <= "11111111";  -- DE4 = FF
      when "0110111100101" =>  data <= "11111111";  -- DE5 = FF
      when "0110111100110" =>  data <= "11111111";  -- DE6 = FF
      when "0110111100111" =>  data <= "11111111";  -- DE7 = FF
      when "0110111101000" =>  data <= "11111111";  -- DE8 = FF
      when "0110111101001" =>  data <= "11111111";  -- DE9 = FF
      when "0110111101010" =>  data <= "11111111";  -- DEA = FF
      when "0110111101011" =>  data <= "11111111";  -- DEB = FF
      when "0110111101100" =>  data <= "11111111";  -- DEC = FF
      when "0110111101101" =>  data <= "11111111";  -- DED = FF
      when "0110111101110" =>  data <= "11111111";  -- DEE = FF
      when "0110111101111" =>  data <= "11111111";  -- DEF = FF
      when "0110111110000" =>  data <= "11111111";  -- DF0 = FF
      when "0110111110001" =>  data <= "11111111";  -- DF1 = FF
      when "0110111110010" =>  data <= "11111111";  -- DF2 = FF
      when "0110111110011" =>  data <= "11111111";  -- DF3 = FF
      when "0110111110100" =>  data <= "11111111";  -- DF4 = FF
      when "0110111110101" =>  data <= "11111111";  -- DF5 = FF
      when "0110111110110" =>  data <= "11111111";  -- DF6 = FF
      when "0110111110111" =>  data <= "11111111";  -- DF7 = FF
      when "0110111111000" =>  data <= "11111111";  -- DF8 = FF
      when "0110111111001" =>  data <= "11111111";  -- DF9 = FF
      when "0110111111010" =>  data <= "11111111";  -- DFA = FF
      when "0110111111011" =>  data <= "11111111";  -- DFB = FF
      when "0110111111100" =>  data <= "11111111";  -- DFC = FF
      when "0110111111101" =>  data <= "11111111";  -- DFD = FF
      when "0110111111110" =>  data <= "11111111";  -- DFE = FF
      when "0110111111111" =>  data <= "11111111";  -- DFF = FF
      when "0111000000000" =>  data <= "11111111";  -- E00 = FF
      when "0111000000001" =>  data <= "11111111";  -- E01 = FF
      when "0111000000010" =>  data <= "11111111";  -- E02 = FF
      when "0111000000011" =>  data <= "11111111";  -- E03 = FF
      when "0111000000100" =>  data <= "11111111";  -- E04 = FF
      when "0111000000101" =>  data <= "11111111";  -- E05 = FF
      when "0111000000110" =>  data <= "11111111";  -- E06 = FF
      when "0111000000111" =>  data <= "11111111";  -- E07 = FF
      when "0111000001000" =>  data <= "11111111";  -- E08 = FF
      when "0111000001001" =>  data <= "11111111";  -- E09 = FF
      when "0111000001010" =>  data <= "11111111";  -- E0A = FF
      when "0111000001011" =>  data <= "11111111";  -- E0B = FF
      when "0111000001100" =>  data <= "11111111";  -- E0C = FF
      when "0111000001101" =>  data <= "11111111";  -- E0D = FF
      when "0111000001110" =>  data <= "11111111";  -- E0E = FF
      when "0111000001111" =>  data <= "11111111";  -- E0F = FF
      when "0111000010000" =>  data <= "11111111";  -- E10 = FF
      when "0111000010001" =>  data <= "11111111";  -- E11 = FF
      when "0111000010010" =>  data <= "11111111";  -- E12 = FF
      when "0111000010011" =>  data <= "11111111";  -- E13 = FF
      when "0111000010100" =>  data <= "11111111";  -- E14 = FF
      when "0111000010101" =>  data <= "11111111";  -- E15 = FF
      when "0111000010110" =>  data <= "11111111";  -- E16 = FF
      when "0111000010111" =>  data <= "11111111";  -- E17 = FF
      when "0111000011000" =>  data <= "11111111";  -- E18 = FF
      when "0111000011001" =>  data <= "11111111";  -- E19 = FF
      when "0111000011010" =>  data <= "11111111";  -- E1A = FF
      when "0111000011011" =>  data <= "11111111";  -- E1B = FF
      when "0111000011100" =>  data <= "11111111";  -- E1C = FF
      when "0111000011101" =>  data <= "11111111";  -- E1D = FF
      when "0111000011110" =>  data <= "11111111";  -- E1E = FF
      when "0111000011111" =>  data <= "11111111";  -- E1F = FF
      when "0111000100000" =>  data <= "11111111";  -- E20 = FF
      when "0111000100001" =>  data <= "11111111";  -- E21 = FF
      when "0111000100010" =>  data <= "11111111";  -- E22 = FF
      when "0111000100011" =>  data <= "11111111";  -- E23 = FF
      when "0111000100100" =>  data <= "11111111";  -- E24 = FF
      when "0111000100101" =>  data <= "11111111";  -- E25 = FF
      when "0111000100110" =>  data <= "11111111";  -- E26 = FF
      when "0111000100111" =>  data <= "11111111";  -- E27 = FF
      when "0111000101000" =>  data <= "11111111";  -- E28 = FF
      when "0111000101001" =>  data <= "11111111";  -- E29 = FF
      when "0111000101010" =>  data <= "11111111";  -- E2A = FF
      when "0111000101011" =>  data <= "11111111";  -- E2B = FF
      when "0111000101100" =>  data <= "11111111";  -- E2C = FF
      when "0111000101101" =>  data <= "11111111";  -- E2D = FF
      when "0111000101110" =>  data <= "11111111";  -- E2E = FF
      when "0111000101111" =>  data <= "11111111";  -- E2F = FF
      when "0111000110000" =>  data <= "11111111";  -- E30 = FF
      when "0111000110001" =>  data <= "11111111";  -- E31 = FF
      when "0111000110010" =>  data <= "11111111";  -- E32 = FF
      when "0111000110011" =>  data <= "11111111";  -- E33 = FF
      when "0111000110100" =>  data <= "11111111";  -- E34 = FF
      when "0111000110101" =>  data <= "11111111";  -- E35 = FF
      when "0111000110110" =>  data <= "11111111";  -- E36 = FF
      when "0111000110111" =>  data <= "11111111";  -- E37 = FF
      when "0111000111000" =>  data <= "11111111";  -- E38 = FF
      when "0111000111001" =>  data <= "11111111";  -- E39 = FF
      when "0111000111010" =>  data <= "11111111";  -- E3A = FF
      when "0111000111011" =>  data <= "11111111";  -- E3B = FF
      when "0111000111100" =>  data <= "11111111";  -- E3C = FF
      when "0111000111101" =>  data <= "11111111";  -- E3D = FF
      when "0111000111110" =>  data <= "11111111";  -- E3E = FF
      when "0111000111111" =>  data <= "11111111";  -- E3F = FF
      when "0111001000000" =>  data <= "11111111";  -- E40 = FF
      when "0111001000001" =>  data <= "11111111";  -- E41 = FF
      when "0111001000010" =>  data <= "11111111";  -- E42 = FF
      when "0111001000011" =>  data <= "11111111";  -- E43 = FF
      when "0111001000100" =>  data <= "11111111";  -- E44 = FF
      when "0111001000101" =>  data <= "11111111";  -- E45 = FF
      when "0111001000110" =>  data <= "11111111";  -- E46 = FF
      when "0111001000111" =>  data <= "11111111";  -- E47 = FF
      when "0111001001000" =>  data <= "11111111";  -- E48 = FF
      when "0111001001001" =>  data <= "11111111";  -- E49 = FF
      when "0111001001010" =>  data <= "11111111";  -- E4A = FF
      when "0111001001011" =>  data <= "11111111";  -- E4B = FF
      when "0111001001100" =>  data <= "11111111";  -- E4C = FF
      when "0111001001101" =>  data <= "11111111";  -- E4D = FF
      when "0111001001110" =>  data <= "11111111";  -- E4E = FF
      when "0111001001111" =>  data <= "11111111";  -- E4F = FF
      when "0111001010000" =>  data <= "11111111";  -- E50 = FF
      when "0111001010001" =>  data <= "11111111";  -- E51 = FF
      when "0111001010010" =>  data <= "11111111";  -- E52 = FF
      when "0111001010011" =>  data <= "11111111";  -- E53 = FF
      when "0111001010100" =>  data <= "11111111";  -- E54 = FF
      when "0111001010101" =>  data <= "11111111";  -- E55 = FF
      when "0111001010110" =>  data <= "11111111";  -- E56 = FF
      when "0111001010111" =>  data <= "11111111";  -- E57 = FF
      when "0111001011000" =>  data <= "11111111";  -- E58 = FF
      when "0111001011001" =>  data <= "11111111";  -- E59 = FF
      when "0111001011010" =>  data <= "11111111";  -- E5A = FF
      when "0111001011011" =>  data <= "11111111";  -- E5B = FF
      when "0111001011100" =>  data <= "11111111";  -- E5C = FF
      when "0111001011101" =>  data <= "11111111";  -- E5D = FF
      when "0111001011110" =>  data <= "11111111";  -- E5E = FF
      when "0111001011111" =>  data <= "11111111";  -- E5F = FF
      when "0111001100000" =>  data <= "11111111";  -- E60 = FF
      when "0111001100001" =>  data <= "11111111";  -- E61 = FF
      when "0111001100010" =>  data <= "11111111";  -- E62 = FF
      when "0111001100011" =>  data <= "11111111";  -- E63 = FF
      when "0111001100100" =>  data <= "11111111";  -- E64 = FF
      when "0111001100101" =>  data <= "11111111";  -- E65 = FF
      when "0111001100110" =>  data <= "11111111";  -- E66 = FF
      when "0111001100111" =>  data <= "11111111";  -- E67 = FF
      when "0111001101000" =>  data <= "11111111";  -- E68 = FF
      when "0111001101001" =>  data <= "11111111";  -- E69 = FF
      when "0111001101010" =>  data <= "11111111";  -- E6A = FF
      when "0111001101011" =>  data <= "11111111";  -- E6B = FF
      when "0111001101100" =>  data <= "11111111";  -- E6C = FF
      when "0111001101101" =>  data <= "11111111";  -- E6D = FF
      when "0111001101110" =>  data <= "11111111";  -- E6E = FF
      when "0111001101111" =>  data <= "11111111";  -- E6F = FF
      when "0111001110000" =>  data <= "11111111";  -- E70 = FF
      when "0111001110001" =>  data <= "11111111";  -- E71 = FF
      when "0111001110010" =>  data <= "11111111";  -- E72 = FF
      when "0111001110011" =>  data <= "11111111";  -- E73 = FF
      when "0111001110100" =>  data <= "11111111";  -- E74 = FF
      when "0111001110101" =>  data <= "11111111";  -- E75 = FF
      when "0111001110110" =>  data <= "11111111";  -- E76 = FF
      when "0111001110111" =>  data <= "11111111";  -- E77 = FF
      when "0111001111000" =>  data <= "11111111";  -- E78 = FF
      when "0111001111001" =>  data <= "11111111";  -- E79 = FF
      when "0111001111010" =>  data <= "11111111";  -- E7A = FF
      when "0111001111011" =>  data <= "11111111";  -- E7B = FF
      when "0111001111100" =>  data <= "11111111";  -- E7C = FF
      when "0111001111101" =>  data <= "11111111";  -- E7D = FF
      when "0111001111110" =>  data <= "11111111";  -- E7E = FF
      when "0111001111111" =>  data <= "11111111";  -- E7F = FF
      when "0111010000000" =>  data <= "11111111";  -- E80 = FF
      when "0111010000001" =>  data <= "11111111";  -- E81 = FF
      when "0111010000010" =>  data <= "11111111";  -- E82 = FF
      when "0111010000011" =>  data <= "11111111";  -- E83 = FF
      when "0111010000100" =>  data <= "11111111";  -- E84 = FF
      when "0111010000101" =>  data <= "11111111";  -- E85 = FF
      when "0111010000110" =>  data <= "11111111";  -- E86 = FF
      when "0111010000111" =>  data <= "11111111";  -- E87 = FF
      when "0111010001000" =>  data <= "11111111";  -- E88 = FF
      when "0111010001001" =>  data <= "11111111";  -- E89 = FF
      when "0111010001010" =>  data <= "11111111";  -- E8A = FF
      when "0111010001011" =>  data <= "11111111";  -- E8B = FF
      when "0111010001100" =>  data <= "11111111";  -- E8C = FF
      when "0111010001101" =>  data <= "11111111";  -- E8D = FF
      when "0111010001110" =>  data <= "11111111";  -- E8E = FF
      when "0111010001111" =>  data <= "11111111";  -- E8F = FF
      when "0111010010000" =>  data <= "11111111";  -- E90 = FF
      when "0111010010001" =>  data <= "11111111";  -- E91 = FF
      when "0111010010010" =>  data <= "11111111";  -- E92 = FF
      when "0111010010011" =>  data <= "11111111";  -- E93 = FF
      when "0111010010100" =>  data <= "11111111";  -- E94 = FF
      when "0111010010101" =>  data <= "11111111";  -- E95 = FF
      when "0111010010110" =>  data <= "11111111";  -- E96 = FF
      when "0111010010111" =>  data <= "11111111";  -- E97 = FF
      when "0111010011000" =>  data <= "11111111";  -- E98 = FF
      when "0111010011001" =>  data <= "11111111";  -- E99 = FF
      when "0111010011010" =>  data <= "11111111";  -- E9A = FF
      when "0111010011011" =>  data <= "11111111";  -- E9B = FF
      when "0111010011100" =>  data <= "11111111";  -- E9C = FF
      when "0111010011101" =>  data <= "11111111";  -- E9D = FF
      when "0111010011110" =>  data <= "11111111";  -- E9E = FF
      when "0111010011111" =>  data <= "11111111";  -- E9F = FF
      when "0111010100000" =>  data <= "11111111";  -- EA0 = FF
      when "0111010100001" =>  data <= "11111111";  -- EA1 = FF
      when "0111010100010" =>  data <= "11111111";  -- EA2 = FF
      when "0111010100011" =>  data <= "11111111";  -- EA3 = FF
      when "0111010100100" =>  data <= "11111111";  -- EA4 = FF
      when "0111010100101" =>  data <= "11111111";  -- EA5 = FF
      when "0111010100110" =>  data <= "11111111";  -- EA6 = FF
      when "0111010100111" =>  data <= "11111111";  -- EA7 = FF
      when "0111010101000" =>  data <= "11111111";  -- EA8 = FF
      when "0111010101001" =>  data <= "11111111";  -- EA9 = FF
      when "0111010101010" =>  data <= "11111111";  -- EAA = FF
      when "0111010101011" =>  data <= "11111111";  -- EAB = FF
      when "0111010101100" =>  data <= "11111111";  -- EAC = FF
      when "0111010101101" =>  data <= "11111111";  -- EAD = FF
      when "0111010101110" =>  data <= "11111111";  -- EAE = FF
      when "0111010101111" =>  data <= "11111111";  -- EAF = FF
      when "0111010110000" =>  data <= "11111111";  -- EB0 = FF
      when "0111010110001" =>  data <= "11111111";  -- EB1 = FF
      when "0111010110010" =>  data <= "11111111";  -- EB2 = FF
      when "0111010110011" =>  data <= "11111111";  -- EB3 = FF
      when "0111010110100" =>  data <= "11111111";  -- EB4 = FF
      when "0111010110101" =>  data <= "11111111";  -- EB5 = FF
      when "0111010110110" =>  data <= "11111111";  -- EB6 = FF
      when "0111010110111" =>  data <= "11111111";  -- EB7 = FF
      when "0111010111000" =>  data <= "11111111";  -- EB8 = FF
      when "0111010111001" =>  data <= "11111111";  -- EB9 = FF
      when "0111010111010" =>  data <= "11111111";  -- EBA = FF
      when "0111010111011" =>  data <= "11111111";  -- EBB = FF
      when "0111010111100" =>  data <= "11111111";  -- EBC = FF
      when "0111010111101" =>  data <= "11111111";  -- EBD = FF
      when "0111010111110" =>  data <= "11111111";  -- EBE = FF
      when "0111010111111" =>  data <= "11111111";  -- EBF = FF
      when "0111011000000" =>  data <= "11111111";  -- EC0 = FF
      when "0111011000001" =>  data <= "11111111";  -- EC1 = FF
      when "0111011000010" =>  data <= "11111111";  -- EC2 = FF
      when "0111011000011" =>  data <= "11111111";  -- EC3 = FF
      when "0111011000100" =>  data <= "11111111";  -- EC4 = FF
      when "0111011000101" =>  data <= "11111111";  -- EC5 = FF
      when "0111011000110" =>  data <= "11111111";  -- EC6 = FF
      when "0111011000111" =>  data <= "11111111";  -- EC7 = FF
      when "0111011001000" =>  data <= "11111111";  -- EC8 = FF
      when "0111011001001" =>  data <= "11111111";  -- EC9 = FF
      when "0111011001010" =>  data <= "11111111";  -- ECA = FF
      when "0111011001011" =>  data <= "11111111";  -- ECB = FF
      when "0111011001100" =>  data <= "11111111";  -- ECC = FF
      when "0111011001101" =>  data <= "11111111";  -- ECD = FF
      when "0111011001110" =>  data <= "11111111";  -- ECE = FF
      when "0111011001111" =>  data <= "11111111";  -- ECF = FF
      when "0111011010000" =>  data <= "11111111";  -- ED0 = FF
      when "0111011010001" =>  data <= "11111111";  -- ED1 = FF
      when "0111011010010" =>  data <= "11111111";  -- ED2 = FF
      when "0111011010011" =>  data <= "11111111";  -- ED3 = FF
      when "0111011010100" =>  data <= "11111111";  -- ED4 = FF
      when "0111011010101" =>  data <= "11111111";  -- ED5 = FF
      when "0111011010110" =>  data <= "11111111";  -- ED6 = FF
      when "0111011010111" =>  data <= "11111111";  -- ED7 = FF
      when "0111011011000" =>  data <= "11111111";  -- ED8 = FF
      when "0111011011001" =>  data <= "11111111";  -- ED9 = FF
      when "0111011011010" =>  data <= "11111111";  -- EDA = FF
      when "0111011011011" =>  data <= "11111111";  -- EDB = FF
      when "0111011011100" =>  data <= "11111111";  -- EDC = FF
      when "0111011011101" =>  data <= "11111111";  -- EDD = FF
      when "0111011011110" =>  data <= "11111111";  -- EDE = FF
      when "0111011011111" =>  data <= "11111111";  -- EDF = FF
      when "0111011100000" =>  data <= "11111111";  -- EE0 = FF
      when "0111011100001" =>  data <= "11111111";  -- EE1 = FF
      when "0111011100010" =>  data <= "11111111";  -- EE2 = FF
      when "0111011100011" =>  data <= "11111111";  -- EE3 = FF
      when "0111011100100" =>  data <= "11111111";  -- EE4 = FF
      when "0111011100101" =>  data <= "11111111";  -- EE5 = FF
      when "0111011100110" =>  data <= "11111111";  -- EE6 = FF
      when "0111011100111" =>  data <= "11111111";  -- EE7 = FF
      when "0111011101000" =>  data <= "11111111";  -- EE8 = FF
      when "0111011101001" =>  data <= "11111111";  -- EE9 = FF
      when "0111011101010" =>  data <= "11111111";  -- EEA = FF
      when "0111011101011" =>  data <= "11111111";  -- EEB = FF
      when "0111011101100" =>  data <= "11111111";  -- EEC = FF
      when "0111011101101" =>  data <= "11111111";  -- EED = FF
      when "0111011101110" =>  data <= "11111111";  -- EEE = FF
      when "0111011101111" =>  data <= "11111111";  -- EEF = FF
      when "0111011110000" =>  data <= "11111111";  -- EF0 = FF
      when "0111011110001" =>  data <= "11111111";  -- EF1 = FF
      when "0111011110010" =>  data <= "11111111";  -- EF2 = FF
      when "0111011110011" =>  data <= "11111111";  -- EF3 = FF
      when "0111011110100" =>  data <= "11111111";  -- EF4 = FF
      when "0111011110101" =>  data <= "11111111";  -- EF5 = FF
      when "0111011110110" =>  data <= "11111111";  -- EF6 = FF
      when "0111011110111" =>  data <= "11111111";  -- EF7 = FF
      when "0111011111000" =>  data <= "11111111";  -- EF8 = FF
      when "0111011111001" =>  data <= "11111111";  -- EF9 = FF
      when "0111011111010" =>  data <= "11111111";  -- EFA = FF
      when "0111011111011" =>  data <= "11111111";  -- EFB = FF
      when "0111011111100" =>  data <= "11111111";  -- EFC = FF
      when "0111011111101" =>  data <= "11111111";  -- EFD = FF
      when "0111011111110" =>  data <= "11111111";  -- EFE = FF
      when "0111011111111" =>  data <= "11111111";  -- EFF = FF
      when "0111100000000" =>  data <= "11111111";  -- F00 = FF
      when "0111100000001" =>  data <= "11111111";  -- F01 = FF
      when "0111100000010" =>  data <= "11111111";  -- F02 = FF
      when "0111100000011" =>  data <= "11111111";  -- F03 = FF
      when "0111100000100" =>  data <= "11111111";  -- F04 = FF
      when "0111100000101" =>  data <= "11111111";  -- F05 = FF
      when "0111100000110" =>  data <= "11111111";  -- F06 = FF
      when "0111100000111" =>  data <= "11111111";  -- F07 = FF
      when "0111100001000" =>  data <= "11111111";  -- F08 = FF
      when "0111100001001" =>  data <= "11111111";  -- F09 = FF
      when "0111100001010" =>  data <= "11111111";  -- F0A = FF
      when "0111100001011" =>  data <= "11111111";  -- F0B = FF
      when "0111100001100" =>  data <= "11111111";  -- F0C = FF
      when "0111100001101" =>  data <= "11111111";  -- F0D = FF
      when "0111100001110" =>  data <= "11111111";  -- F0E = FF
      when "0111100001111" =>  data <= "11111111";  -- F0F = FF
      when "0111100010000" =>  data <= "11111111";  -- F10 = FF
      when "0111100010001" =>  data <= "11111111";  -- F11 = FF
      when "0111100010010" =>  data <= "11111111";  -- F12 = FF
      when "0111100010011" =>  data <= "11111111";  -- F13 = FF
      when "0111100010100" =>  data <= "11111111";  -- F14 = FF
      when "0111100010101" =>  data <= "11111111";  -- F15 = FF
      when "0111100010110" =>  data <= "11111111";  -- F16 = FF
      when "0111100010111" =>  data <= "11111111";  -- F17 = FF
      when "0111100011000" =>  data <= "11111111";  -- F18 = FF
      when "0111100011001" =>  data <= "11111111";  -- F19 = FF
      when "0111100011010" =>  data <= "11111111";  -- F1A = FF
      when "0111100011011" =>  data <= "11111111";  -- F1B = FF
      when "0111100011100" =>  data <= "11111111";  -- F1C = FF
      when "0111100011101" =>  data <= "11111111";  -- F1D = FF
      when "0111100011110" =>  data <= "11111111";  -- F1E = FF
      when "0111100011111" =>  data <= "11111111";  -- F1F = FF
      when "0111100100000" =>  data <= "11111111";  -- F20 = FF
      when "0111100100001" =>  data <= "11111111";  -- F21 = FF
      when "0111100100010" =>  data <= "11111111";  -- F22 = FF
      when "0111100100011" =>  data <= "11111111";  -- F23 = FF
      when "0111100100100" =>  data <= "11111111";  -- F24 = FF
      when "0111100100101" =>  data <= "11111111";  -- F25 = FF
      when "0111100100110" =>  data <= "11111111";  -- F26 = FF
      when "0111100100111" =>  data <= "11111111";  -- F27 = FF
      when "0111100101000" =>  data <= "11111111";  -- F28 = FF
      when "0111100101001" =>  data <= "11111111";  -- F29 = FF
      when "0111100101010" =>  data <= "11111111";  -- F2A = FF
      when "0111100101011" =>  data <= "11111111";  -- F2B = FF
      when "0111100101100" =>  data <= "11111111";  -- F2C = FF
      when "0111100101101" =>  data <= "11111111";  -- F2D = FF
      when "0111100101110" =>  data <= "11111111";  -- F2E = FF
      when "0111100101111" =>  data <= "11111111";  -- F2F = FF
      when "0111100110000" =>  data <= "11111111";  -- F30 = FF
      when "0111100110001" =>  data <= "11111111";  -- F31 = FF
      when "0111100110010" =>  data <= "11111111";  -- F32 = FF
      when "0111100110011" =>  data <= "11111111";  -- F33 = FF
      when "0111100110100" =>  data <= "11111111";  -- F34 = FF
      when "0111100110101" =>  data <= "11111111";  -- F35 = FF
      when "0111100110110" =>  data <= "11111111";  -- F36 = FF
      when "0111100110111" =>  data <= "11111111";  -- F37 = FF
      when "0111100111000" =>  data <= "11111111";  -- F38 = FF
      when "0111100111001" =>  data <= "11111111";  -- F39 = FF
      when "0111100111010" =>  data <= "11111111";  -- F3A = FF
      when "0111100111011" =>  data <= "11111111";  -- F3B = FF
      when "0111100111100" =>  data <= "11111111";  -- F3C = FF
      when "0111100111101" =>  data <= "11111111";  -- F3D = FF
      when "0111100111110" =>  data <= "11111111";  -- F3E = FF
      when "0111100111111" =>  data <= "11111111";  -- F3F = FF
      when "0111101000000" =>  data <= "11111111";  -- F40 = FF
      when "0111101000001" =>  data <= "11111111";  -- F41 = FF
      when "0111101000010" =>  data <= "11111111";  -- F42 = FF
      when "0111101000011" =>  data <= "11111111";  -- F43 = FF
      when "0111101000100" =>  data <= "11111111";  -- F44 = FF
      when "0111101000101" =>  data <= "11111111";  -- F45 = FF
      when "0111101000110" =>  data <= "11111111";  -- F46 = FF
      when "0111101000111" =>  data <= "11111111";  -- F47 = FF
      when "0111101001000" =>  data <= "11111111";  -- F48 = FF
      when "0111101001001" =>  data <= "11111111";  -- F49 = FF
      when "0111101001010" =>  data <= "11111111";  -- F4A = FF
      when "0111101001011" =>  data <= "11111111";  -- F4B = FF
      when "0111101001100" =>  data <= "11111111";  -- F4C = FF
      when "0111101001101" =>  data <= "11111111";  -- F4D = FF
      when "0111101001110" =>  data <= "11111111";  -- F4E = FF
      when "0111101001111" =>  data <= "11111111";  -- F4F = FF
      when "0111101010000" =>  data <= "11111111";  -- F50 = FF
      when "0111101010001" =>  data <= "11111111";  -- F51 = FF
      when "0111101010010" =>  data <= "11111111";  -- F52 = FF
      when "0111101010011" =>  data <= "11111111";  -- F53 = FF
      when "0111101010100" =>  data <= "11111111";  -- F54 = FF
      when "0111101010101" =>  data <= "11111111";  -- F55 = FF
      when "0111101010110" =>  data <= "11111111";  -- F56 = FF
      when "0111101010111" =>  data <= "11111111";  -- F57 = FF
      when "0111101011000" =>  data <= "11111111";  -- F58 = FF
      when "0111101011001" =>  data <= "11111111";  -- F59 = FF
      when "0111101011010" =>  data <= "11111111";  -- F5A = FF
      when "0111101011011" =>  data <= "11111111";  -- F5B = FF
      when "0111101011100" =>  data <= "11111111";  -- F5C = FF
      when "0111101011101" =>  data <= "11111111";  -- F5D = FF
      when "0111101011110" =>  data <= "11111111";  -- F5E = FF
      when "0111101011111" =>  data <= "11111111";  -- F5F = FF
      when "0111101100000" =>  data <= "11111111";  -- F60 = FF
      when "0111101100001" =>  data <= "11111111";  -- F61 = FF
      when "0111101100010" =>  data <= "11111111";  -- F62 = FF
      when "0111101100011" =>  data <= "11111111";  -- F63 = FF
      when "0111101100100" =>  data <= "11111111";  -- F64 = FF
      when "0111101100101" =>  data <= "11111111";  -- F65 = FF
      when "0111101100110" =>  data <= "11111111";  -- F66 = FF
      when "0111101100111" =>  data <= "11111111";  -- F67 = FF
      when "0111101101000" =>  data <= "11111111";  -- F68 = FF
      when "0111101101001" =>  data <= "11111111";  -- F69 = FF
      when "0111101101010" =>  data <= "11111111";  -- F6A = FF
      when "0111101101011" =>  data <= "11111111";  -- F6B = FF
      when "0111101101100" =>  data <= "11111111";  -- F6C = FF
      when "0111101101101" =>  data <= "11111111";  -- F6D = FF
      when "0111101101110" =>  data <= "11111111";  -- F6E = FF
      when "0111101101111" =>  data <= "11111111";  -- F6F = FF
      when "0111101110000" =>  data <= "11111111";  -- F70 = FF
      when "0111101110001" =>  data <= "11111111";  -- F71 = FF
      when "0111101110010" =>  data <= "11111111";  -- F72 = FF
      when "0111101110011" =>  data <= "11111111";  -- F73 = FF
      when "0111101110100" =>  data <= "11111111";  -- F74 = FF
      when "0111101110101" =>  data <= "11111111";  -- F75 = FF
      when "0111101110110" =>  data <= "11111111";  -- F76 = FF
      when "0111101110111" =>  data <= "11111111";  -- F77 = FF
      when "0111101111000" =>  data <= "11111111";  -- F78 = FF
      when "0111101111001" =>  data <= "11111111";  -- F79 = FF
      when "0111101111010" =>  data <= "11111111";  -- F7A = FF
      when "0111101111011" =>  data <= "11111111";  -- F7B = FF
      when "0111101111100" =>  data <= "11111111";  -- F7C = FF
      when "0111101111101" =>  data <= "11111111";  -- F7D = FF
      when "0111101111110" =>  data <= "11111111";  -- F7E = FF
      when "0111101111111" =>  data <= "11111111";  -- F7F = FF
      when "0111110000000" =>  data <= "11111111";  -- F80 = FF
      when "0111110000001" =>  data <= "11111111";  -- F81 = FF
      when "0111110000010" =>  data <= "11111111";  -- F82 = FF
      when "0111110000011" =>  data <= "11111111";  -- F83 = FF
      when "0111110000100" =>  data <= "11111111";  -- F84 = FF
      when "0111110000101" =>  data <= "11111111";  -- F85 = FF
      when "0111110000110" =>  data <= "11111111";  -- F86 = FF
      when "0111110000111" =>  data <= "11111111";  -- F87 = FF
      when "0111110001000" =>  data <= "11111111";  -- F88 = FF
      when "0111110001001" =>  data <= "11111111";  -- F89 = FF
      when "0111110001010" =>  data <= "11111111";  -- F8A = FF
      when "0111110001011" =>  data <= "11111111";  -- F8B = FF
      when "0111110001100" =>  data <= "11111111";  -- F8C = FF
      when "0111110001101" =>  data <= "11111111";  -- F8D = FF
      when "0111110001110" =>  data <= "11111111";  -- F8E = FF
      when "0111110001111" =>  data <= "11111111";  -- F8F = FF
      when "0111110010000" =>  data <= "11111111";  -- F90 = FF
      when "0111110010001" =>  data <= "11111111";  -- F91 = FF
      when "0111110010010" =>  data <= "11111111";  -- F92 = FF
      when "0111110010011" =>  data <= "11111111";  -- F93 = FF
      when "0111110010100" =>  data <= "11111111";  -- F94 = FF
      when "0111110010101" =>  data <= "11111111";  -- F95 = FF
      when "0111110010110" =>  data <= "11111111";  -- F96 = FF
      when "0111110010111" =>  data <= "11111111";  -- F97 = FF
      when "0111110011000" =>  data <= "11111111";  -- F98 = FF
      when "0111110011001" =>  data <= "11111111";  -- F99 = FF
      when "0111110011010" =>  data <= "11111111";  -- F9A = FF
      when "0111110011011" =>  data <= "11111111";  -- F9B = FF
      when "0111110011100" =>  data <= "11111111";  -- F9C = FF
      when "0111110011101" =>  data <= "11111111";  -- F9D = FF
      when "0111110011110" =>  data <= "11111111";  -- F9E = FF
      when "0111110011111" =>  data <= "11111111";  -- F9F = FF
      when "0111110100000" =>  data <= "11111111";  -- FA0 = FF
      when "0111110100001" =>  data <= "11111111";  -- FA1 = FF
      when "0111110100010" =>  data <= "11111111";  -- FA2 = FF
      when "0111110100011" =>  data <= "11111111";  -- FA3 = FF
      when "0111110100100" =>  data <= "11111111";  -- FA4 = FF
      when "0111110100101" =>  data <= "11111111";  -- FA5 = FF
      when "0111110100110" =>  data <= "11111111";  -- FA6 = FF
      when "0111110100111" =>  data <= "11111111";  -- FA7 = FF
      when "0111110101000" =>  data <= "11111111";  -- FA8 = FF
      when "0111110101001" =>  data <= "11111111";  -- FA9 = FF
      when "0111110101010" =>  data <= "11111111";  -- FAA = FF
      when "0111110101011" =>  data <= "11111111";  -- FAB = FF
      when "0111110101100" =>  data <= "11111111";  -- FAC = FF
      when "0111110101101" =>  data <= "11111111";  -- FAD = FF
      when "0111110101110" =>  data <= "11111111";  -- FAE = FF
      when "0111110101111" =>  data <= "11111111";  -- FAF = FF
      when "0111110110000" =>  data <= "11111111";  -- FB0 = FF
      when "0111110110001" =>  data <= "11111111";  -- FB1 = FF
      when "0111110110010" =>  data <= "11111111";  -- FB2 = FF
      when "0111110110011" =>  data <= "11111111";  -- FB3 = FF
      when "0111110110100" =>  data <= "11111111";  -- FB4 = FF
      when "0111110110101" =>  data <= "11111111";  -- FB5 = FF
      when "0111110110110" =>  data <= "11111111";  -- FB6 = FF
      when "0111110110111" =>  data <= "11111111";  -- FB7 = FF
      when "0111110111000" =>  data <= "11111111";  -- FB8 = FF
      when "0111110111001" =>  data <= "11111111";  -- FB9 = FF
      when "0111110111010" =>  data <= "11111111";  -- FBA = FF
      when "0111110111011" =>  data <= "11111111";  -- FBB = FF
      when "0111110111100" =>  data <= "11111111";  -- FBC = FF
      when "0111110111101" =>  data <= "11111111";  -- FBD = FF
      when "0111110111110" =>  data <= "11111111";  -- FBE = FF
      when "0111110111111" =>  data <= "11111111";  -- FBF = FF
      when "0111111000000" =>  data <= "11111111";  -- FC0 = FF
      when "0111111000001" =>  data <= "11111111";  -- FC1 = FF
      when "0111111000010" =>  data <= "11111111";  -- FC2 = FF
      when "0111111000011" =>  data <= "11111111";  -- FC3 = FF
      when "0111111000100" =>  data <= "11111111";  -- FC4 = FF
      when "0111111000101" =>  data <= "11111111";  -- FC5 = FF
      when "0111111000110" =>  data <= "11111111";  -- FC6 = FF
      when "0111111000111" =>  data <= "11111111";  -- FC7 = FF
      when "0111111001000" =>  data <= "11111111";  -- FC8 = FF
      when "0111111001001" =>  data <= "11111111";  -- FC9 = FF
      when "0111111001010" =>  data <= "11111111";  -- FCA = FF
      when "0111111001011" =>  data <= "11111111";  -- FCB = FF
      when "0111111001100" =>  data <= "11111111";  -- FCC = FF
      when "0111111001101" =>  data <= "11111111";  -- FCD = FF
      when "0111111001110" =>  data <= "11111111";  -- FCE = FF
      when "0111111001111" =>  data <= "11111111";  -- FCF = FF
      when "0111111010000" =>  data <= "11111111";  -- FD0 = FF
      when "0111111010001" =>  data <= "11111111";  -- FD1 = FF
      when "0111111010010" =>  data <= "11111111";  -- FD2 = FF
      when "0111111010011" =>  data <= "11111111";  -- FD3 = FF
      when "0111111010100" =>  data <= "11111111";  -- FD4 = FF
      when "0111111010101" =>  data <= "11111111";  -- FD5 = FF
      when "0111111010110" =>  data <= "11111111";  -- FD6 = FF
      when "0111111010111" =>  data <= "11111111";  -- FD7 = FF
      when "0111111011000" =>  data <= "11111111";  -- FD8 = FF
      when "0111111011001" =>  data <= "11111111";  -- FD9 = FF
      when "0111111011010" =>  data <= "11111111";  -- FDA = FF
      when "0111111011011" =>  data <= "11111111";  -- FDB = FF
      when "0111111011100" =>  data <= "11111111";  -- FDC = FF
      when "0111111011101" =>  data <= "11111111";  -- FDD = FF
      when "0111111011110" =>  data <= "11111111";  -- FDE = FF
      when "0111111011111" =>  data <= "11111111";  -- FDF = FF
      when "0111111100000" =>  data <= "11111111";  -- FE0 = FF
      when "0111111100001" =>  data <= "11111111";  -- FE1 = FF
      when "0111111100010" =>  data <= "11111111";  -- FE2 = FF
      when "0111111100011" =>  data <= "11111111";  -- FE3 = FF
      when "0111111100100" =>  data <= "11111111";  -- FE4 = FF
      when "0111111100101" =>  data <= "11111111";  -- FE5 = FF
      when "0111111100110" =>  data <= "11111111";  -- FE6 = FF
      when "0111111100111" =>  data <= "11111111";  -- FE7 = FF
      when "0111111101000" =>  data <= "11111111";  -- FE8 = FF
      when "0111111101001" =>  data <= "11111111";  -- FE9 = FF
      when "0111111101010" =>  data <= "11111111";  -- FEA = FF
      when "0111111101011" =>  data <= "11111111";  -- FEB = FF
      when "0111111101100" =>  data <= "11111111";  -- FEC = FF
      when "0111111101101" =>  data <= "11111111";  -- FED = FF
      when "0111111101110" =>  data <= "11111111";  -- FEE = FF
      when "0111111101111" =>  data <= "11111111";  -- FEF = FF
      when "0111111110000" =>  data <= "11111111";  -- FF0 = FF
      when "0111111110001" =>  data <= "11111111";  -- FF1 = FF
      when "0111111110010" =>  data <= "11111111";  -- FF2 = FF
      when "0111111110011" =>  data <= "11111111";  -- FF3 = FF
      when "0111111110100" =>  data <= "11111111";  -- FF4 = FF
      when "0111111110101" =>  data <= "11111111";  -- FF5 = FF
      when "0111111110110" =>  data <= "11111111";  -- FF6 = FF
      when "0111111110111" =>  data <= "11111111";  -- FF7 = FF
      when "0111111111000" =>  data <= "11111111";  -- FF8 = FF
      when "0111111111001" =>  data <= "11111111";  -- FF9 = FF
      when "0111111111010" =>  data <= "11111111";  -- FFA = FF
      when "0111111111011" =>  data <= "11111111";  -- FFB = FF
      when "0111111111100" =>  data <= "11111111";  -- FFC = FF
      when "0111111111101" =>  data <= "11111111";  -- FFD = FF
      when "0111111111110" =>  data <= "11111111";  -- FFE = FF
      when "0111111111111" =>  data <= "11111111";  -- FFF = FF
      when "1000000000000" =>  data <= "11111111";  -- 1000 = FF
      when "1000000000001" =>  data <= "11111111";  -- 1001 = FF
      when "1000000000010" =>  data <= "11111111";  -- 1002 = FF
      when "1000000000011" =>  data <= "11111111";  -- 1003 = FF
      when "1000000000100" =>  data <= "11111111";  -- 1004 = FF
      when "1000000000101" =>  data <= "11111111";  -- 1005 = FF
      when "1000000000110" =>  data <= "11111111";  -- 1006 = FF
      when "1000000000111" =>  data <= "11111111";  -- 1007 = FF
      when "1000000001000" =>  data <= "11111111";  -- 1008 = FF
      when "1000000001001" =>  data <= "11111111";  -- 1009 = FF
      when "1000000001010" =>  data <= "11111111";  -- 100A = FF
      when "1000000001011" =>  data <= "11111111";  -- 100B = FF
      when "1000000001100" =>  data <= "11111111";  -- 100C = FF
      when "1000000001101" =>  data <= "11111111";  -- 100D = FF
      when "1000000001110" =>  data <= "11111111";  -- 100E = FF
      when "1000000001111" =>  data <= "11111111";  -- 100F = FF
      when "1000000010000" =>  data <= "11111111";  -- 1010 = FF
      when "1000000010001" =>  data <= "11111111";  -- 1011 = FF
      when "1000000010010" =>  data <= "11111111";  -- 1012 = FF
      when "1000000010011" =>  data <= "11111111";  -- 1013 = FF
      when "1000000010100" =>  data <= "11111111";  -- 1014 = FF
      when "1000000010101" =>  data <= "11111111";  -- 1015 = FF
      when "1000000010110" =>  data <= "11111111";  -- 1016 = FF
      when "1000000010111" =>  data <= "11111111";  -- 1017 = FF
      when "1000000011000" =>  data <= "11111111";  -- 1018 = FF
      when "1000000011001" =>  data <= "11111111";  -- 1019 = FF
      when "1000000011010" =>  data <= "11111111";  -- 101A = FF
      when "1000000011011" =>  data <= "11111111";  -- 101B = FF
      when "1000000011100" =>  data <= "11111111";  -- 101C = FF
      when "1000000011101" =>  data <= "11111111";  -- 101D = FF
      when "1000000011110" =>  data <= "11111111";  -- 101E = FF
      when "1000000011111" =>  data <= "11111111";  -- 101F = FF
      when "1000000100000" =>  data <= "11111111";  -- 1020 = FF
      when "1000000100001" =>  data <= "11111111";  -- 1021 = FF
      when "1000000100010" =>  data <= "11111111";  -- 1022 = FF
      when "1000000100011" =>  data <= "11111111";  -- 1023 = FF
      when "1000000100100" =>  data <= "11111111";  -- 1024 = FF
      when "1000000100101" =>  data <= "11111111";  -- 1025 = FF
      when "1000000100110" =>  data <= "11111111";  -- 1026 = FF
      when "1000000100111" =>  data <= "11111111";  -- 1027 = FF
      when "1000000101000" =>  data <= "11111111";  -- 1028 = FF
      when "1000000101001" =>  data <= "11111111";  -- 1029 = FF
      when "1000000101010" =>  data <= "11111111";  -- 102A = FF
      when "1000000101011" =>  data <= "11111111";  -- 102B = FF
      when "1000000101100" =>  data <= "11111111";  -- 102C = FF
      when "1000000101101" =>  data <= "11111111";  -- 102D = FF
      when "1000000101110" =>  data <= "11111111";  -- 102E = FF
      when "1000000101111" =>  data <= "11111111";  -- 102F = FF
      when "1000000110000" =>  data <= "11111111";  -- 1030 = FF
      when "1000000110001" =>  data <= "11111111";  -- 1031 = FF
      when "1000000110010" =>  data <= "11111111";  -- 1032 = FF
      when "1000000110011" =>  data <= "11111111";  -- 1033 = FF
      when "1000000110100" =>  data <= "11111111";  -- 1034 = FF
      when "1000000110101" =>  data <= "11111111";  -- 1035 = FF
      when "1000000110110" =>  data <= "11111111";  -- 1036 = FF
      when "1000000110111" =>  data <= "11111111";  -- 1037 = FF
      when "1000000111000" =>  data <= "11111111";  -- 1038 = FF
      when "1000000111001" =>  data <= "11111111";  -- 1039 = FF
      when "1000000111010" =>  data <= "11111111";  -- 103A = FF
      when "1000000111011" =>  data <= "11111111";  -- 103B = FF
      when "1000000111100" =>  data <= "11111111";  -- 103C = FF
      when "1000000111101" =>  data <= "11111111";  -- 103D = FF
      when "1000000111110" =>  data <= "11111111";  -- 103E = FF
      when "1000000111111" =>  data <= "11111111";  -- 103F = FF
      when "1000001000000" =>  data <= "11111111";  -- 1040 = FF
      when "1000001000001" =>  data <= "11111111";  -- 1041 = FF
      when "1000001000010" =>  data <= "11111111";  -- 1042 = FF
      when "1000001000011" =>  data <= "11111111";  -- 1043 = FF
      when "1000001000100" =>  data <= "11111111";  -- 1044 = FF
      when "1000001000101" =>  data <= "11111111";  -- 1045 = FF
      when "1000001000110" =>  data <= "11111111";  -- 1046 = FF
      when "1000001000111" =>  data <= "11111111";  -- 1047 = FF
      when "1000001001000" =>  data <= "11111111";  -- 1048 = FF
      when "1000001001001" =>  data <= "11111111";  -- 1049 = FF
      when "1000001001010" =>  data <= "11111111";  -- 104A = FF
      when "1000001001011" =>  data <= "11111111";  -- 104B = FF
      when "1000001001100" =>  data <= "11111111";  -- 104C = FF
      when "1000001001101" =>  data <= "11111111";  -- 104D = FF
      when "1000001001110" =>  data <= "11111111";  -- 104E = FF
      when "1000001001111" =>  data <= "11111111";  -- 104F = FF
      when "1000001010000" =>  data <= "11111111";  -- 1050 = FF
      when "1000001010001" =>  data <= "11111111";  -- 1051 = FF
      when "1000001010010" =>  data <= "11111111";  -- 1052 = FF
      when "1000001010011" =>  data <= "11111111";  -- 1053 = FF
      when "1000001010100" =>  data <= "11111111";  -- 1054 = FF
      when "1000001010101" =>  data <= "11111111";  -- 1055 = FF
      when "1000001010110" =>  data <= "11111111";  -- 1056 = FF
      when "1000001010111" =>  data <= "11111111";  -- 1057 = FF
      when "1000001011000" =>  data <= "11111111";  -- 1058 = FF
      when "1000001011001" =>  data <= "11111111";  -- 1059 = FF
      when "1000001011010" =>  data <= "11111111";  -- 105A = FF
      when "1000001011011" =>  data <= "11111111";  -- 105B = FF
      when "1000001011100" =>  data <= "11111111";  -- 105C = FF
      when "1000001011101" =>  data <= "11111111";  -- 105D = FF
      when "1000001011110" =>  data <= "11111111";  -- 105E = FF
      when "1000001011111" =>  data <= "11111111";  -- 105F = FF
      when "1000001100000" =>  data <= "11111111";  -- 1060 = FF
      when "1000001100001" =>  data <= "11111111";  -- 1061 = FF
      when "1000001100010" =>  data <= "11111111";  -- 1062 = FF
      when "1000001100011" =>  data <= "11111111";  -- 1063 = FF
      when "1000001100100" =>  data <= "11111111";  -- 1064 = FF
      when "1000001100101" =>  data <= "11111111";  -- 1065 = FF
      when "1000001100110" =>  data <= "11111111";  -- 1066 = FF
      when "1000001100111" =>  data <= "11111111";  -- 1067 = FF
      when "1000001101000" =>  data <= "11111111";  -- 1068 = FF
      when "1000001101001" =>  data <= "11111111";  -- 1069 = FF
      when "1000001101010" =>  data <= "11111111";  -- 106A = FF
      when "1000001101011" =>  data <= "11111111";  -- 106B = FF
      when "1000001101100" =>  data <= "11111111";  -- 106C = FF
      when "1000001101101" =>  data <= "11111111";  -- 106D = FF
      when "1000001101110" =>  data <= "11111111";  -- 106E = FF
      when "1000001101111" =>  data <= "11111111";  -- 106F = FF
      when "1000001110000" =>  data <= "11111111";  -- 1070 = FF
      when "1000001110001" =>  data <= "11111111";  -- 1071 = FF
      when "1000001110010" =>  data <= "11111111";  -- 1072 = FF
      when "1000001110011" =>  data <= "11111111";  -- 1073 = FF
      when "1000001110100" =>  data <= "11111111";  -- 1074 = FF
      when "1000001110101" =>  data <= "11111111";  -- 1075 = FF
      when "1000001110110" =>  data <= "11111111";  -- 1076 = FF
      when "1000001110111" =>  data <= "11111111";  -- 1077 = FF
      when "1000001111000" =>  data <= "11111111";  -- 1078 = FF
      when "1000001111001" =>  data <= "11111111";  -- 1079 = FF
      when "1000001111010" =>  data <= "11111111";  -- 107A = FF
      when "1000001111011" =>  data <= "11111111";  -- 107B = FF
      when "1000001111100" =>  data <= "11111111";  -- 107C = FF
      when "1000001111101" =>  data <= "11111111";  -- 107D = FF
      when "1000001111110" =>  data <= "11111111";  -- 107E = FF
      when "1000001111111" =>  data <= "11111111";  -- 107F = FF
      when "1000010000000" =>  data <= "11111111";  -- 1080 = FF
      when "1000010000001" =>  data <= "11111111";  -- 1081 = FF
      when "1000010000010" =>  data <= "11111111";  -- 1082 = FF
      when "1000010000011" =>  data <= "11111111";  -- 1083 = FF
      when "1000010000100" =>  data <= "11111111";  -- 1084 = FF
      when "1000010000101" =>  data <= "11111111";  -- 1085 = FF
      when "1000010000110" =>  data <= "11111111";  -- 1086 = FF
      when "1000010000111" =>  data <= "11111111";  -- 1087 = FF
      when "1000010001000" =>  data <= "11111111";  -- 1088 = FF
      when "1000010001001" =>  data <= "11111111";  -- 1089 = FF
      when "1000010001010" =>  data <= "11111111";  -- 108A = FF
      when "1000010001011" =>  data <= "11111111";  -- 108B = FF
      when "1000010001100" =>  data <= "11111111";  -- 108C = FF
      when "1000010001101" =>  data <= "11111111";  -- 108D = FF
      when "1000010001110" =>  data <= "11111111";  -- 108E = FF
      when "1000010001111" =>  data <= "11111111";  -- 108F = FF
      when "1000010010000" =>  data <= "11111111";  -- 1090 = FF
      when "1000010010001" =>  data <= "11111111";  -- 1091 = FF
      when "1000010010010" =>  data <= "11111111";  -- 1092 = FF
      when "1000010010011" =>  data <= "11111111";  -- 1093 = FF
      when "1000010010100" =>  data <= "11111111";  -- 1094 = FF
      when "1000010010101" =>  data <= "11111111";  -- 1095 = FF
      when "1000010010110" =>  data <= "11111111";  -- 1096 = FF
      when "1000010010111" =>  data <= "11111111";  -- 1097 = FF
      when "1000010011000" =>  data <= "11111111";  -- 1098 = FF
      when "1000010011001" =>  data <= "11111111";  -- 1099 = FF
      when "1000010011010" =>  data <= "11111111";  -- 109A = FF
      when "1000010011011" =>  data <= "11111111";  -- 109B = FF
      when "1000010011100" =>  data <= "11111111";  -- 109C = FF
      when "1000010011101" =>  data <= "11111111";  -- 109D = FF
      when "1000010011110" =>  data <= "11111111";  -- 109E = FF
      when "1000010011111" =>  data <= "11111111";  -- 109F = FF
      when "1000010100000" =>  data <= "11111111";  -- 10A0 = FF
      when "1000010100001" =>  data <= "11111111";  -- 10A1 = FF
      when "1000010100010" =>  data <= "11111111";  -- 10A2 = FF
      when "1000010100011" =>  data <= "11111111";  -- 10A3 = FF
      when "1000010100100" =>  data <= "11111111";  -- 10A4 = FF
      when "1000010100101" =>  data <= "11111111";  -- 10A5 = FF
      when "1000010100110" =>  data <= "11111111";  -- 10A6 = FF
      when "1000010100111" =>  data <= "11111111";  -- 10A7 = FF
      when "1000010101000" =>  data <= "11111111";  -- 10A8 = FF
      when "1000010101001" =>  data <= "11111111";  -- 10A9 = FF
      when "1000010101010" =>  data <= "11111111";  -- 10AA = FF
      when "1000010101011" =>  data <= "11111111";  -- 10AB = FF
      when "1000010101100" =>  data <= "11111111";  -- 10AC = FF
      when "1000010101101" =>  data <= "11111111";  -- 10AD = FF
      when "1000010101110" =>  data <= "11111111";  -- 10AE = FF
      when "1000010101111" =>  data <= "11111111";  -- 10AF = FF
      when "1000010110000" =>  data <= "11111111";  -- 10B0 = FF
      when "1000010110001" =>  data <= "11111111";  -- 10B1 = FF
      when "1000010110010" =>  data <= "11111111";  -- 10B2 = FF
      when "1000010110011" =>  data <= "11111111";  -- 10B3 = FF
      when "1000010110100" =>  data <= "11111111";  -- 10B4 = FF
      when "1000010110101" =>  data <= "11111111";  -- 10B5 = FF
      when "1000010110110" =>  data <= "11111111";  -- 10B6 = FF
      when "1000010110111" =>  data <= "11111111";  -- 10B7 = FF
      when "1000010111000" =>  data <= "11111111";  -- 10B8 = FF
      when "1000010111001" =>  data <= "11111111";  -- 10B9 = FF
      when "1000010111010" =>  data <= "11111111";  -- 10BA = FF
      when "1000010111011" =>  data <= "11111111";  -- 10BB = FF
      when "1000010111100" =>  data <= "11111111";  -- 10BC = FF
      when "1000010111101" =>  data <= "11111111";  -- 10BD = FF
      when "1000010111110" =>  data <= "11111111";  -- 10BE = FF
      when "1000010111111" =>  data <= "11111111";  -- 10BF = FF
      when "1000011000000" =>  data <= "11111111";  -- 10C0 = FF
      when "1000011000001" =>  data <= "11111111";  -- 10C1 = FF
      when "1000011000010" =>  data <= "11111111";  -- 10C2 = FF
      when "1000011000011" =>  data <= "11111111";  -- 10C3 = FF
      when "1000011000100" =>  data <= "11111111";  -- 10C4 = FF
      when "1000011000101" =>  data <= "11111111";  -- 10C5 = FF
      when "1000011000110" =>  data <= "11111111";  -- 10C6 = FF
      when "1000011000111" =>  data <= "11111111";  -- 10C7 = FF
      when "1000011001000" =>  data <= "11111111";  -- 10C8 = FF
      when "1000011001001" =>  data <= "11111111";  -- 10C9 = FF
      when "1000011001010" =>  data <= "11111111";  -- 10CA = FF
      when "1000011001011" =>  data <= "11111111";  -- 10CB = FF
      when "1000011001100" =>  data <= "11111111";  -- 10CC = FF
      when "1000011001101" =>  data <= "11111111";  -- 10CD = FF
      when "1000011001110" =>  data <= "11111111";  -- 10CE = FF
      when "1000011001111" =>  data <= "11111111";  -- 10CF = FF
      when "1000011010000" =>  data <= "11111111";  -- 10D0 = FF
      when "1000011010001" =>  data <= "11111111";  -- 10D1 = FF
      when "1000011010010" =>  data <= "11111111";  -- 10D2 = FF
      when "1000011010011" =>  data <= "11111111";  -- 10D3 = FF
      when "1000011010100" =>  data <= "11111111";  -- 10D4 = FF
      when "1000011010101" =>  data <= "11111111";  -- 10D5 = FF
      when "1000011010110" =>  data <= "11111111";  -- 10D6 = FF
      when "1000011010111" =>  data <= "11111111";  -- 10D7 = FF
      when "1000011011000" =>  data <= "11111111";  -- 10D8 = FF
      when "1000011011001" =>  data <= "11111111";  -- 10D9 = FF
      when "1000011011010" =>  data <= "11111111";  -- 10DA = FF
      when "1000011011011" =>  data <= "11111111";  -- 10DB = FF
      when "1000011011100" =>  data <= "11111111";  -- 10DC = FF
      when "1000011011101" =>  data <= "11111111";  -- 10DD = FF
      when "1000011011110" =>  data <= "11111111";  -- 10DE = FF
      when "1000011011111" =>  data <= "11111111";  -- 10DF = FF
      when "1000011100000" =>  data <= "11111111";  -- 10E0 = FF
      when "1000011100001" =>  data <= "11111111";  -- 10E1 = FF
      when "1000011100010" =>  data <= "11111111";  -- 10E2 = FF
      when "1000011100011" =>  data <= "11111111";  -- 10E3 = FF
      when "1000011100100" =>  data <= "11111111";  -- 10E4 = FF
      when "1000011100101" =>  data <= "11111111";  -- 10E5 = FF
      when "1000011100110" =>  data <= "11111111";  -- 10E6 = FF
      when "1000011100111" =>  data <= "11111111";  -- 10E7 = FF
      when "1000011101000" =>  data <= "11111111";  -- 10E8 = FF
      when "1000011101001" =>  data <= "11111111";  -- 10E9 = FF
      when "1000011101010" =>  data <= "11111111";  -- 10EA = FF
      when "1000011101011" =>  data <= "11111111";  -- 10EB = FF
      when "1000011101100" =>  data <= "11111111";  -- 10EC = FF
      when "1000011101101" =>  data <= "11111111";  -- 10ED = FF
      when "1000011101110" =>  data <= "11111111";  -- 10EE = FF
      when "1000011101111" =>  data <= "11111111";  -- 10EF = FF
      when "1000011110000" =>  data <= "11111111";  -- 10F0 = FF
      when "1000011110001" =>  data <= "11111111";  -- 10F1 = FF
      when "1000011110010" =>  data <= "11111111";  -- 10F2 = FF
      when "1000011110011" =>  data <= "11111111";  -- 10F3 = FF
      when "1000011110100" =>  data <= "11111111";  -- 10F4 = FF
      when "1000011110101" =>  data <= "11111111";  -- 10F5 = FF
      when "1000011110110" =>  data <= "11111111";  -- 10F6 = FF
      when "1000011110111" =>  data <= "11111111";  -- 10F7 = FF
      when "1000011111000" =>  data <= "11111111";  -- 10F8 = FF
      when "1000011111001" =>  data <= "11111111";  -- 10F9 = FF
      when "1000011111010" =>  data <= "11111111";  -- 10FA = FF
      when "1000011111011" =>  data <= "11111111";  -- 10FB = FF
      when "1000011111100" =>  data <= "11111111";  -- 10FC = FF
      when "1000011111101" =>  data <= "11111111";  -- 10FD = FF
      when "1000011111110" =>  data <= "11111111";  -- 10FE = FF
      when "1000011111111" =>  data <= "11111111";  -- 10FF = FF
      when "1000100000000" =>  data <= "11111111";  -- 1100 = FF
      when "1000100000001" =>  data <= "11111111";  -- 1101 = FF
      when "1000100000010" =>  data <= "11111111";  -- 1102 = FF
      when "1000100000011" =>  data <= "11111111";  -- 1103 = FF
      when "1000100000100" =>  data <= "11111111";  -- 1104 = FF
      when "1000100000101" =>  data <= "11111111";  -- 1105 = FF
      when "1000100000110" =>  data <= "11111111";  -- 1106 = FF
      when "1000100000111" =>  data <= "11111111";  -- 1107 = FF
      when "1000100001000" =>  data <= "11111111";  -- 1108 = FF
      when "1000100001001" =>  data <= "11111111";  -- 1109 = FF
      when "1000100001010" =>  data <= "11111111";  -- 110A = FF
      when "1000100001011" =>  data <= "11111111";  -- 110B = FF
      when "1000100001100" =>  data <= "11111111";  -- 110C = FF
      when "1000100001101" =>  data <= "11111111";  -- 110D = FF
      when "1000100001110" =>  data <= "11111111";  -- 110E = FF
      when "1000100001111" =>  data <= "11111111";  -- 110F = FF
      when "1000100010000" =>  data <= "11111111";  -- 1110 = FF
      when "1000100010001" =>  data <= "11111111";  -- 1111 = FF
      when "1000100010010" =>  data <= "11111111";  -- 1112 = FF
      when "1000100010011" =>  data <= "11111111";  -- 1113 = FF
      when "1000100010100" =>  data <= "11111111";  -- 1114 = FF
      when "1000100010101" =>  data <= "11111111";  -- 1115 = FF
      when "1000100010110" =>  data <= "11111111";  -- 1116 = FF
      when "1000100010111" =>  data <= "11111111";  -- 1117 = FF
      when "1000100011000" =>  data <= "11111111";  -- 1118 = FF
      when "1000100011001" =>  data <= "11111111";  -- 1119 = FF
      when "1000100011010" =>  data <= "11111111";  -- 111A = FF
      when "1000100011011" =>  data <= "11111111";  -- 111B = FF
      when "1000100011100" =>  data <= "11111111";  -- 111C = FF
      when "1000100011101" =>  data <= "11111111";  -- 111D = FF
      when "1000100011110" =>  data <= "11111111";  -- 111E = FF
      when "1000100011111" =>  data <= "11111111";  -- 111F = FF
      when "1000100100000" =>  data <= "11111111";  -- 1120 = FF
      when "1000100100001" =>  data <= "11111111";  -- 1121 = FF
      when "1000100100010" =>  data <= "11111111";  -- 1122 = FF
      when "1000100100011" =>  data <= "11111111";  -- 1123 = FF
      when "1000100100100" =>  data <= "11111111";  -- 1124 = FF
      when "1000100100101" =>  data <= "11111111";  -- 1125 = FF
      when "1000100100110" =>  data <= "11111111";  -- 1126 = FF
      when "1000100100111" =>  data <= "11111111";  -- 1127 = FF
      when "1000100101000" =>  data <= "11111111";  -- 1128 = FF
      when "1000100101001" =>  data <= "11111111";  -- 1129 = FF
      when "1000100101010" =>  data <= "11111111";  -- 112A = FF
      when "1000100101011" =>  data <= "11111111";  -- 112B = FF
      when "1000100101100" =>  data <= "11111111";  -- 112C = FF
      when "1000100101101" =>  data <= "11111111";  -- 112D = FF
      when "1000100101110" =>  data <= "11111111";  -- 112E = FF
      when "1000100101111" =>  data <= "11111111";  -- 112F = FF
      when "1000100110000" =>  data <= "11111111";  -- 1130 = FF
      when "1000100110001" =>  data <= "11111111";  -- 1131 = FF
      when "1000100110010" =>  data <= "11111111";  -- 1132 = FF
      when "1000100110011" =>  data <= "11111111";  -- 1133 = FF
      when "1000100110100" =>  data <= "11111111";  -- 1134 = FF
      when "1000100110101" =>  data <= "11111111";  -- 1135 = FF
      when "1000100110110" =>  data <= "11111111";  -- 1136 = FF
      when "1000100110111" =>  data <= "11111111";  -- 1137 = FF
      when "1000100111000" =>  data <= "11111111";  -- 1138 = FF
      when "1000100111001" =>  data <= "11111111";  -- 1139 = FF
      when "1000100111010" =>  data <= "11111111";  -- 113A = FF
      when "1000100111011" =>  data <= "11111111";  -- 113B = FF
      when "1000100111100" =>  data <= "11111111";  -- 113C = FF
      when "1000100111101" =>  data <= "11111111";  -- 113D = FF
      when "1000100111110" =>  data <= "11111111";  -- 113E = FF
      when "1000100111111" =>  data <= "11111111";  -- 113F = FF
      when "1000101000000" =>  data <= "11111111";  -- 1140 = FF
      when "1000101000001" =>  data <= "11111111";  -- 1141 = FF
      when "1000101000010" =>  data <= "11111111";  -- 1142 = FF
      when "1000101000011" =>  data <= "11111111";  -- 1143 = FF
      when "1000101000100" =>  data <= "11111111";  -- 1144 = FF
      when "1000101000101" =>  data <= "11111111";  -- 1145 = FF
      when "1000101000110" =>  data <= "11111111";  -- 1146 = FF
      when "1000101000111" =>  data <= "11111111";  -- 1147 = FF
      when "1000101001000" =>  data <= "11111111";  -- 1148 = FF
      when "1000101001001" =>  data <= "11111111";  -- 1149 = FF
      when "1000101001010" =>  data <= "11111111";  -- 114A = FF
      when "1000101001011" =>  data <= "11111111";  -- 114B = FF
      when "1000101001100" =>  data <= "11111111";  -- 114C = FF
      when "1000101001101" =>  data <= "11111111";  -- 114D = FF
      when "1000101001110" =>  data <= "11111111";  -- 114E = FF
      when "1000101001111" =>  data <= "11111111";  -- 114F = FF
      when "1000101010000" =>  data <= "11111111";  -- 1150 = FF
      when "1000101010001" =>  data <= "11111111";  -- 1151 = FF
      when "1000101010010" =>  data <= "11111111";  -- 1152 = FF
      when "1000101010011" =>  data <= "11111111";  -- 1153 = FF
      when "1000101010100" =>  data <= "11111111";  -- 1154 = FF
      when "1000101010101" =>  data <= "11111111";  -- 1155 = FF
      when "1000101010110" =>  data <= "11111111";  -- 1156 = FF
      when "1000101010111" =>  data <= "11111111";  -- 1157 = FF
      when "1000101011000" =>  data <= "11111111";  -- 1158 = FF
      when "1000101011001" =>  data <= "11111111";  -- 1159 = FF
      when "1000101011010" =>  data <= "11111111";  -- 115A = FF
      when "1000101011011" =>  data <= "11111111";  -- 115B = FF
      when "1000101011100" =>  data <= "11111111";  -- 115C = FF
      when "1000101011101" =>  data <= "11111111";  -- 115D = FF
      when "1000101011110" =>  data <= "11111111";  -- 115E = FF
      when "1000101011111" =>  data <= "11111111";  -- 115F = FF
      when "1000101100000" =>  data <= "11111111";  -- 1160 = FF
      when "1000101100001" =>  data <= "11111111";  -- 1161 = FF
      when "1000101100010" =>  data <= "11111111";  -- 1162 = FF
      when "1000101100011" =>  data <= "11111111";  -- 1163 = FF
      when "1000101100100" =>  data <= "11111111";  -- 1164 = FF
      when "1000101100101" =>  data <= "11111111";  -- 1165 = FF
      when "1000101100110" =>  data <= "11111111";  -- 1166 = FF
      when "1000101100111" =>  data <= "11111111";  -- 1167 = FF
      when "1000101101000" =>  data <= "11111111";  -- 1168 = FF
      when "1000101101001" =>  data <= "11111111";  -- 1169 = FF
      when "1000101101010" =>  data <= "11111111";  -- 116A = FF
      when "1000101101011" =>  data <= "11111111";  -- 116B = FF
      when "1000101101100" =>  data <= "11111111";  -- 116C = FF
      when "1000101101101" =>  data <= "11111111";  -- 116D = FF
      when "1000101101110" =>  data <= "11111111";  -- 116E = FF
      when "1000101101111" =>  data <= "11111111";  -- 116F = FF
      when "1000101110000" =>  data <= "11111111";  -- 1170 = FF
      when "1000101110001" =>  data <= "11111111";  -- 1171 = FF
      when "1000101110010" =>  data <= "11111111";  -- 1172 = FF
      when "1000101110011" =>  data <= "11111111";  -- 1173 = FF
      when "1000101110100" =>  data <= "11111111";  -- 1174 = FF
      when "1000101110101" =>  data <= "11111111";  -- 1175 = FF
      when "1000101110110" =>  data <= "11111111";  -- 1176 = FF
      when "1000101110111" =>  data <= "11111111";  -- 1177 = FF
      when "1000101111000" =>  data <= "11111111";  -- 1178 = FF
      when "1000101111001" =>  data <= "11111111";  -- 1179 = FF
      when "1000101111010" =>  data <= "11111111";  -- 117A = FF
      when "1000101111011" =>  data <= "11111111";  -- 117B = FF
      when "1000101111100" =>  data <= "11111111";  -- 117C = FF
      when "1000101111101" =>  data <= "11111111";  -- 117D = FF
      when "1000101111110" =>  data <= "11111111";  -- 117E = FF
      when "1000101111111" =>  data <= "11111111";  -- 117F = FF
      when "1000110000000" =>  data <= "11111111";  -- 1180 = FF
      when "1000110000001" =>  data <= "11111111";  -- 1181 = FF
      when "1000110000010" =>  data <= "11111111";  -- 1182 = FF
      when "1000110000011" =>  data <= "11111111";  -- 1183 = FF
      when "1000110000100" =>  data <= "11111111";  -- 1184 = FF
      when "1000110000101" =>  data <= "11111111";  -- 1185 = FF
      when "1000110000110" =>  data <= "11111111";  -- 1186 = FF
      when "1000110000111" =>  data <= "11111111";  -- 1187 = FF
      when "1000110001000" =>  data <= "11111111";  -- 1188 = FF
      when "1000110001001" =>  data <= "11111111";  -- 1189 = FF
      when "1000110001010" =>  data <= "11111111";  -- 118A = FF
      when "1000110001011" =>  data <= "11111111";  -- 118B = FF
      when "1000110001100" =>  data <= "11111111";  -- 118C = FF
      when "1000110001101" =>  data <= "11111111";  -- 118D = FF
      when "1000110001110" =>  data <= "11111111";  -- 118E = FF
      when "1000110001111" =>  data <= "11111111";  -- 118F = FF
      when "1000110010000" =>  data <= "11111111";  -- 1190 = FF
      when "1000110010001" =>  data <= "11111111";  -- 1191 = FF
      when "1000110010010" =>  data <= "11111111";  -- 1192 = FF
      when "1000110010011" =>  data <= "11111111";  -- 1193 = FF
      when "1000110010100" =>  data <= "11111111";  -- 1194 = FF
      when "1000110010101" =>  data <= "11111111";  -- 1195 = FF
      when "1000110010110" =>  data <= "11111111";  -- 1196 = FF
      when "1000110010111" =>  data <= "11111111";  -- 1197 = FF
      when "1000110011000" =>  data <= "11111111";  -- 1198 = FF
      when "1000110011001" =>  data <= "11111111";  -- 1199 = FF
      when "1000110011010" =>  data <= "11111111";  -- 119A = FF
      when "1000110011011" =>  data <= "11111111";  -- 119B = FF
      when "1000110011100" =>  data <= "11111111";  -- 119C = FF
      when "1000110011101" =>  data <= "11111111";  -- 119D = FF
      when "1000110011110" =>  data <= "11111111";  -- 119E = FF
      when "1000110011111" =>  data <= "11111111";  -- 119F = FF
      when "1000110100000" =>  data <= "11111111";  -- 11A0 = FF
      when "1000110100001" =>  data <= "11111111";  -- 11A1 = FF
      when "1000110100010" =>  data <= "11111111";  -- 11A2 = FF
      when "1000110100011" =>  data <= "11111111";  -- 11A3 = FF
      when "1000110100100" =>  data <= "11111111";  -- 11A4 = FF
      when "1000110100101" =>  data <= "11111111";  -- 11A5 = FF
      when "1000110100110" =>  data <= "11111111";  -- 11A6 = FF
      when "1000110100111" =>  data <= "11111111";  -- 11A7 = FF
      when "1000110101000" =>  data <= "11111111";  -- 11A8 = FF
      when "1000110101001" =>  data <= "11111111";  -- 11A9 = FF
      when "1000110101010" =>  data <= "11111111";  -- 11AA = FF
      when "1000110101011" =>  data <= "11111111";  -- 11AB = FF
      when "1000110101100" =>  data <= "11111111";  -- 11AC = FF
      when "1000110101101" =>  data <= "11111111";  -- 11AD = FF
      when "1000110101110" =>  data <= "11111111";  -- 11AE = FF
      when "1000110101111" =>  data <= "11111111";  -- 11AF = FF
      when "1000110110000" =>  data <= "11111111";  -- 11B0 = FF
      when "1000110110001" =>  data <= "11111111";  -- 11B1 = FF
      when "1000110110010" =>  data <= "11111111";  -- 11B2 = FF
      when "1000110110011" =>  data <= "11111111";  -- 11B3 = FF
      when "1000110110100" =>  data <= "11111111";  -- 11B4 = FF
      when "1000110110101" =>  data <= "11111111";  -- 11B5 = FF
      when "1000110110110" =>  data <= "11111111";  -- 11B6 = FF
      when "1000110110111" =>  data <= "11111111";  -- 11B7 = FF
      when "1000110111000" =>  data <= "11111111";  -- 11B8 = FF
      when "1000110111001" =>  data <= "11111111";  -- 11B9 = FF
      when "1000110111010" =>  data <= "11111111";  -- 11BA = FF
      when "1000110111011" =>  data <= "11111111";  -- 11BB = FF
      when "1000110111100" =>  data <= "11111111";  -- 11BC = FF
      when "1000110111101" =>  data <= "11111111";  -- 11BD = FF
      when "1000110111110" =>  data <= "11111111";  -- 11BE = FF
      when "1000110111111" =>  data <= "11111111";  -- 11BF = FF
      when "1000111000000" =>  data <= "11111111";  -- 11C0 = FF
      when "1000111000001" =>  data <= "11111111";  -- 11C1 = FF
      when "1000111000010" =>  data <= "11111111";  -- 11C2 = FF
      when "1000111000011" =>  data <= "11111111";  -- 11C3 = FF
      when "1000111000100" =>  data <= "11111111";  -- 11C4 = FF
      when "1000111000101" =>  data <= "11111111";  -- 11C5 = FF
      when "1000111000110" =>  data <= "11111111";  -- 11C6 = FF
      when "1000111000111" =>  data <= "11111111";  -- 11C7 = FF
      when "1000111001000" =>  data <= "11111111";  -- 11C8 = FF
      when "1000111001001" =>  data <= "11111111";  -- 11C9 = FF
      when "1000111001010" =>  data <= "11111111";  -- 11CA = FF
      when "1000111001011" =>  data <= "11111111";  -- 11CB = FF
      when "1000111001100" =>  data <= "11111111";  -- 11CC = FF
      when "1000111001101" =>  data <= "11111111";  -- 11CD = FF
      when "1000111001110" =>  data <= "11111111";  -- 11CE = FF
      when "1000111001111" =>  data <= "11111111";  -- 11CF = FF
      when "1000111010000" =>  data <= "11111111";  -- 11D0 = FF
      when "1000111010001" =>  data <= "11111111";  -- 11D1 = FF
      when "1000111010010" =>  data <= "11111111";  -- 11D2 = FF
      when "1000111010011" =>  data <= "11111111";  -- 11D3 = FF
      when "1000111010100" =>  data <= "11111111";  -- 11D4 = FF
      when "1000111010101" =>  data <= "11111111";  -- 11D5 = FF
      when "1000111010110" =>  data <= "11111111";  -- 11D6 = FF
      when "1000111010111" =>  data <= "11111111";  -- 11D7 = FF
      when "1000111011000" =>  data <= "11111111";  -- 11D8 = FF
      when "1000111011001" =>  data <= "11111111";  -- 11D9 = FF
      when "1000111011010" =>  data <= "11111111";  -- 11DA = FF
      when "1000111011011" =>  data <= "11111111";  -- 11DB = FF
      when "1000111011100" =>  data <= "11111111";  -- 11DC = FF
      when "1000111011101" =>  data <= "11111111";  -- 11DD = FF
      when "1000111011110" =>  data <= "11111111";  -- 11DE = FF
      when "1000111011111" =>  data <= "11111111";  -- 11DF = FF
      when "1000111100000" =>  data <= "11111111";  -- 11E0 = FF
      when "1000111100001" =>  data <= "11111111";  -- 11E1 = FF
      when "1000111100010" =>  data <= "11111111";  -- 11E2 = FF
      when "1000111100011" =>  data <= "11111111";  -- 11E3 = FF
      when "1000111100100" =>  data <= "11111111";  -- 11E4 = FF
      when "1000111100101" =>  data <= "11111111";  -- 11E5 = FF
      when "1000111100110" =>  data <= "11111111";  -- 11E6 = FF
      when "1000111100111" =>  data <= "11111111";  -- 11E7 = FF
      when "1000111101000" =>  data <= "11111111";  -- 11E8 = FF
      when "1000111101001" =>  data <= "11111111";  -- 11E9 = FF
      when "1000111101010" =>  data <= "11111111";  -- 11EA = FF
      when "1000111101011" =>  data <= "11111111";  -- 11EB = FF
      when "1000111101100" =>  data <= "11111111";  -- 11EC = FF
      when "1000111101101" =>  data <= "11111111";  -- 11ED = FF
      when "1000111101110" =>  data <= "11111111";  -- 11EE = FF
      when "1000111101111" =>  data <= "11111111";  -- 11EF = FF
      when "1000111110000" =>  data <= "11111111";  -- 11F0 = FF
      when "1000111110001" =>  data <= "11111111";  -- 11F1 = FF
      when "1000111110010" =>  data <= "11111111";  -- 11F2 = FF
      when "1000111110011" =>  data <= "11111111";  -- 11F3 = FF
      when "1000111110100" =>  data <= "11111111";  -- 11F4 = FF
      when "1000111110101" =>  data <= "11111111";  -- 11F5 = FF
      when "1000111110110" =>  data <= "11111111";  -- 11F6 = FF
      when "1000111110111" =>  data <= "11111111";  -- 11F7 = FF
      when "1000111111000" =>  data <= "11111111";  -- 11F8 = FF
      when "1000111111001" =>  data <= "11111111";  -- 11F9 = FF
      when "1000111111010" =>  data <= "11111111";  -- 11FA = FF
      when "1000111111011" =>  data <= "11111111";  -- 11FB = FF
      when "1000111111100" =>  data <= "11111111";  -- 11FC = FF
      when "1000111111101" =>  data <= "11111111";  -- 11FD = FF
      when "1000111111110" =>  data <= "11111111";  -- 11FE = FF
      when "1000111111111" =>  data <= "11111111";  -- 11FF = FF
      when "1001000000000" =>  data <= "11111111";  -- 1200 = FF
      when "1001000000001" =>  data <= "11111111";  -- 1201 = FF
      when "1001000000010" =>  data <= "11111111";  -- 1202 = FF
      when "1001000000011" =>  data <= "11111111";  -- 1203 = FF
      when "1001000000100" =>  data <= "11111111";  -- 1204 = FF
      when "1001000000101" =>  data <= "11111111";  -- 1205 = FF
      when "1001000000110" =>  data <= "11111111";  -- 1206 = FF
      when "1001000000111" =>  data <= "11111111";  -- 1207 = FF
      when "1001000001000" =>  data <= "11111111";  -- 1208 = FF
      when "1001000001001" =>  data <= "11111111";  -- 1209 = FF
      when "1001000001010" =>  data <= "11111111";  -- 120A = FF
      when "1001000001011" =>  data <= "11111111";  -- 120B = FF
      when "1001000001100" =>  data <= "11111111";  -- 120C = FF
      when "1001000001101" =>  data <= "11111111";  -- 120D = FF
      when "1001000001110" =>  data <= "11111111";  -- 120E = FF
      when "1001000001111" =>  data <= "11111111";  -- 120F = FF
      when "1001000010000" =>  data <= "11111111";  -- 1210 = FF
      when "1001000010001" =>  data <= "11111111";  -- 1211 = FF
      when "1001000010010" =>  data <= "11111111";  -- 1212 = FF
      when "1001000010011" =>  data <= "11111111";  -- 1213 = FF
      when "1001000010100" =>  data <= "11111111";  -- 1214 = FF
      when "1001000010101" =>  data <= "11111111";  -- 1215 = FF
      when "1001000010110" =>  data <= "11111111";  -- 1216 = FF
      when "1001000010111" =>  data <= "11111111";  -- 1217 = FF
      when "1001000011000" =>  data <= "11111111";  -- 1218 = FF
      when "1001000011001" =>  data <= "11111111";  -- 1219 = FF
      when "1001000011010" =>  data <= "11111111";  -- 121A = FF
      when "1001000011011" =>  data <= "11111111";  -- 121B = FF
      when "1001000011100" =>  data <= "11111111";  -- 121C = FF
      when "1001000011101" =>  data <= "11111111";  -- 121D = FF
      when "1001000011110" =>  data <= "11111111";  -- 121E = FF
      when "1001000011111" =>  data <= "11111111";  -- 121F = FF
      when "1001000100000" =>  data <= "11111111";  -- 1220 = FF
      when "1001000100001" =>  data <= "11111111";  -- 1221 = FF
      when "1001000100010" =>  data <= "11111111";  -- 1222 = FF
      when "1001000100011" =>  data <= "11111111";  -- 1223 = FF
      when "1001000100100" =>  data <= "11111111";  -- 1224 = FF
      when "1001000100101" =>  data <= "11111111";  -- 1225 = FF
      when "1001000100110" =>  data <= "11111111";  -- 1226 = FF
      when "1001000100111" =>  data <= "11111111";  -- 1227 = FF
      when "1001000101000" =>  data <= "11111111";  -- 1228 = FF
      when "1001000101001" =>  data <= "11111111";  -- 1229 = FF
      when "1001000101010" =>  data <= "11111111";  -- 122A = FF
      when "1001000101011" =>  data <= "11111111";  -- 122B = FF
      when "1001000101100" =>  data <= "11111111";  -- 122C = FF
      when "1001000101101" =>  data <= "11111111";  -- 122D = FF
      when "1001000101110" =>  data <= "11111111";  -- 122E = FF
      when "1001000101111" =>  data <= "11111111";  -- 122F = FF
      when "1001000110000" =>  data <= "11111111";  -- 1230 = FF
      when "1001000110001" =>  data <= "11111111";  -- 1231 = FF
      when "1001000110010" =>  data <= "11111111";  -- 1232 = FF
      when "1001000110011" =>  data <= "11111111";  -- 1233 = FF
      when "1001000110100" =>  data <= "11111111";  -- 1234 = FF
      when "1001000110101" =>  data <= "11111111";  -- 1235 = FF
      when "1001000110110" =>  data <= "11111111";  -- 1236 = FF
      when "1001000110111" =>  data <= "11111111";  -- 1237 = FF
      when "1001000111000" =>  data <= "11111111";  -- 1238 = FF
      when "1001000111001" =>  data <= "11111111";  -- 1239 = FF
      when "1001000111010" =>  data <= "11111111";  -- 123A = FF
      when "1001000111011" =>  data <= "11111111";  -- 123B = FF
      when "1001000111100" =>  data <= "11111111";  -- 123C = FF
      when "1001000111101" =>  data <= "11111111";  -- 123D = FF
      when "1001000111110" =>  data <= "11111111";  -- 123E = FF
      when "1001000111111" =>  data <= "11111111";  -- 123F = FF
      when "1001001000000" =>  data <= "11111111";  -- 1240 = FF
      when "1001001000001" =>  data <= "11111111";  -- 1241 = FF
      when "1001001000010" =>  data <= "11111111";  -- 1242 = FF
      when "1001001000011" =>  data <= "11111111";  -- 1243 = FF
      when "1001001000100" =>  data <= "11111111";  -- 1244 = FF
      when "1001001000101" =>  data <= "11111111";  -- 1245 = FF
      when "1001001000110" =>  data <= "11111111";  -- 1246 = FF
      when "1001001000111" =>  data <= "11111111";  -- 1247 = FF
      when "1001001001000" =>  data <= "11111111";  -- 1248 = FF
      when "1001001001001" =>  data <= "11111111";  -- 1249 = FF
      when "1001001001010" =>  data <= "11111111";  -- 124A = FF
      when "1001001001011" =>  data <= "11111111";  -- 124B = FF
      when "1001001001100" =>  data <= "11111111";  -- 124C = FF
      when "1001001001101" =>  data <= "11111111";  -- 124D = FF
      when "1001001001110" =>  data <= "11111111";  -- 124E = FF
      when "1001001001111" =>  data <= "11111111";  -- 124F = FF
      when "1001001010000" =>  data <= "11111111";  -- 1250 = FF
      when "1001001010001" =>  data <= "11111111";  -- 1251 = FF
      when "1001001010010" =>  data <= "11111111";  -- 1252 = FF
      when "1001001010011" =>  data <= "11111111";  -- 1253 = FF
      when "1001001010100" =>  data <= "11111111";  -- 1254 = FF
      when "1001001010101" =>  data <= "11111111";  -- 1255 = FF
      when "1001001010110" =>  data <= "11111111";  -- 1256 = FF
      when "1001001010111" =>  data <= "11111111";  -- 1257 = FF
      when "1001001011000" =>  data <= "11111111";  -- 1258 = FF
      when "1001001011001" =>  data <= "11111111";  -- 1259 = FF
      when "1001001011010" =>  data <= "11111111";  -- 125A = FF
      when "1001001011011" =>  data <= "11111111";  -- 125B = FF
      when "1001001011100" =>  data <= "11111111";  -- 125C = FF
      when "1001001011101" =>  data <= "11111111";  -- 125D = FF
      when "1001001011110" =>  data <= "11111111";  -- 125E = FF
      when "1001001011111" =>  data <= "11111111";  -- 125F = FF
      when "1001001100000" =>  data <= "11111111";  -- 1260 = FF
      when "1001001100001" =>  data <= "11111111";  -- 1261 = FF
      when "1001001100010" =>  data <= "11111111";  -- 1262 = FF
      when "1001001100011" =>  data <= "11111111";  -- 1263 = FF
      when "1001001100100" =>  data <= "11111111";  -- 1264 = FF
      when "1001001100101" =>  data <= "11111111";  -- 1265 = FF
      when "1001001100110" =>  data <= "11111111";  -- 1266 = FF
      when "1001001100111" =>  data <= "11111111";  -- 1267 = FF
      when "1001001101000" =>  data <= "11111111";  -- 1268 = FF
      when "1001001101001" =>  data <= "11111111";  -- 1269 = FF
      when "1001001101010" =>  data <= "11111111";  -- 126A = FF
      when "1001001101011" =>  data <= "11111111";  -- 126B = FF
      when "1001001101100" =>  data <= "11111111";  -- 126C = FF
      when "1001001101101" =>  data <= "11111111";  -- 126D = FF
      when "1001001101110" =>  data <= "11111111";  -- 126E = FF
      when "1001001101111" =>  data <= "11111111";  -- 126F = FF
      when "1001001110000" =>  data <= "11111111";  -- 1270 = FF
      when "1001001110001" =>  data <= "11111111";  -- 1271 = FF
      when "1001001110010" =>  data <= "11111111";  -- 1272 = FF
      when "1001001110011" =>  data <= "11111111";  -- 1273 = FF
      when "1001001110100" =>  data <= "11111111";  -- 1274 = FF
      when "1001001110101" =>  data <= "11111111";  -- 1275 = FF
      when "1001001110110" =>  data <= "11111111";  -- 1276 = FF
      when "1001001110111" =>  data <= "11111111";  -- 1277 = FF
      when "1001001111000" =>  data <= "11111111";  -- 1278 = FF
      when "1001001111001" =>  data <= "11111111";  -- 1279 = FF
      when "1001001111010" =>  data <= "11111111";  -- 127A = FF
      when "1001001111011" =>  data <= "11111111";  -- 127B = FF
      when "1001001111100" =>  data <= "11111111";  -- 127C = FF
      when "1001001111101" =>  data <= "11111111";  -- 127D = FF
      when "1001001111110" =>  data <= "11111111";  -- 127E = FF
      when "1001001111111" =>  data <= "11111111";  -- 127F = FF
      when "1001010000000" =>  data <= "11111111";  -- 1280 = FF
      when "1001010000001" =>  data <= "11111111";  -- 1281 = FF
      when "1001010000010" =>  data <= "11111111";  -- 1282 = FF
      when "1001010000011" =>  data <= "11111111";  -- 1283 = FF
      when "1001010000100" =>  data <= "11111111";  -- 1284 = FF
      when "1001010000101" =>  data <= "11111111";  -- 1285 = FF
      when "1001010000110" =>  data <= "11111111";  -- 1286 = FF
      when "1001010000111" =>  data <= "11111111";  -- 1287 = FF
      when "1001010001000" =>  data <= "11111111";  -- 1288 = FF
      when "1001010001001" =>  data <= "11111111";  -- 1289 = FF
      when "1001010001010" =>  data <= "11111111";  -- 128A = FF
      when "1001010001011" =>  data <= "11111111";  -- 128B = FF
      when "1001010001100" =>  data <= "11111111";  -- 128C = FF
      when "1001010001101" =>  data <= "11111111";  -- 128D = FF
      when "1001010001110" =>  data <= "11111111";  -- 128E = FF
      when "1001010001111" =>  data <= "11111111";  -- 128F = FF
      when "1001010010000" =>  data <= "11111111";  -- 1290 = FF
      when "1001010010001" =>  data <= "11111111";  -- 1291 = FF
      when "1001010010010" =>  data <= "11111111";  -- 1292 = FF
      when "1001010010011" =>  data <= "11111111";  -- 1293 = FF
      when "1001010010100" =>  data <= "11111111";  -- 1294 = FF
      when "1001010010101" =>  data <= "11111111";  -- 1295 = FF
      when "1001010010110" =>  data <= "11111111";  -- 1296 = FF
      when "1001010010111" =>  data <= "11111111";  -- 1297 = FF
      when "1001010011000" =>  data <= "11111111";  -- 1298 = FF
      when "1001010011001" =>  data <= "11111111";  -- 1299 = FF
      when "1001010011010" =>  data <= "11111111";  -- 129A = FF
      when "1001010011011" =>  data <= "11111111";  -- 129B = FF
      when "1001010011100" =>  data <= "11111111";  -- 129C = FF
      when "1001010011101" =>  data <= "11111111";  -- 129D = FF
      when "1001010011110" =>  data <= "11111111";  -- 129E = FF
      when "1001010011111" =>  data <= "11111111";  -- 129F = FF
      when "1001010100000" =>  data <= "11111111";  -- 12A0 = FF
      when "1001010100001" =>  data <= "11111111";  -- 12A1 = FF
      when "1001010100010" =>  data <= "11111111";  -- 12A2 = FF
      when "1001010100011" =>  data <= "11111111";  -- 12A3 = FF
      when "1001010100100" =>  data <= "11111111";  -- 12A4 = FF
      when "1001010100101" =>  data <= "11111111";  -- 12A5 = FF
      when "1001010100110" =>  data <= "11111111";  -- 12A6 = FF
      when "1001010100111" =>  data <= "11111111";  -- 12A7 = FF
      when "1001010101000" =>  data <= "11111111";  -- 12A8 = FF
      when "1001010101001" =>  data <= "11111111";  -- 12A9 = FF
      when "1001010101010" =>  data <= "11111111";  -- 12AA = FF
      when "1001010101011" =>  data <= "11111111";  -- 12AB = FF
      when "1001010101100" =>  data <= "11111111";  -- 12AC = FF
      when "1001010101101" =>  data <= "11111111";  -- 12AD = FF
      when "1001010101110" =>  data <= "11111111";  -- 12AE = FF
      when "1001010101111" =>  data <= "11111111";  -- 12AF = FF
      when "1001010110000" =>  data <= "11111111";  -- 12B0 = FF
      when "1001010110001" =>  data <= "11111111";  -- 12B1 = FF
      when "1001010110010" =>  data <= "11111111";  -- 12B2 = FF
      when "1001010110011" =>  data <= "11111111";  -- 12B3 = FF
      when "1001010110100" =>  data <= "11111111";  -- 12B4 = FF
      when "1001010110101" =>  data <= "11111111";  -- 12B5 = FF
      when "1001010110110" =>  data <= "11111111";  -- 12B6 = FF
      when "1001010110111" =>  data <= "11111111";  -- 12B7 = FF
      when "1001010111000" =>  data <= "11111111";  -- 12B8 = FF
      when "1001010111001" =>  data <= "11111111";  -- 12B9 = FF
      when "1001010111010" =>  data <= "11111111";  -- 12BA = FF
      when "1001010111011" =>  data <= "11111111";  -- 12BB = FF
      when "1001010111100" =>  data <= "11111111";  -- 12BC = FF
      when "1001010111101" =>  data <= "11111111";  -- 12BD = FF
      when "1001010111110" =>  data <= "11111111";  -- 12BE = FF
      when "1001010111111" =>  data <= "11111111";  -- 12BF = FF
      when "1001011000000" =>  data <= "11111111";  -- 12C0 = FF
      when "1001011000001" =>  data <= "11111111";  -- 12C1 = FF
      when "1001011000010" =>  data <= "11111111";  -- 12C2 = FF
      when "1001011000011" =>  data <= "11111111";  -- 12C3 = FF
      when "1001011000100" =>  data <= "11111111";  -- 12C4 = FF
      when "1001011000101" =>  data <= "11111111";  -- 12C5 = FF
      when "1001011000110" =>  data <= "11111111";  -- 12C6 = FF
      when "1001011000111" =>  data <= "11111111";  -- 12C7 = FF
      when "1001011001000" =>  data <= "11111111";  -- 12C8 = FF
      when "1001011001001" =>  data <= "11111111";  -- 12C9 = FF
      when "1001011001010" =>  data <= "11111111";  -- 12CA = FF
      when "1001011001011" =>  data <= "11111111";  -- 12CB = FF
      when "1001011001100" =>  data <= "11111111";  -- 12CC = FF
      when "1001011001101" =>  data <= "11111111";  -- 12CD = FF
      when "1001011001110" =>  data <= "11111111";  -- 12CE = FF
      when "1001011001111" =>  data <= "11111111";  -- 12CF = FF
      when "1001011010000" =>  data <= "11111111";  -- 12D0 = FF
      when "1001011010001" =>  data <= "11111111";  -- 12D1 = FF
      when "1001011010010" =>  data <= "11111111";  -- 12D2 = FF
      when "1001011010011" =>  data <= "11111111";  -- 12D3 = FF
      when "1001011010100" =>  data <= "11111111";  -- 12D4 = FF
      when "1001011010101" =>  data <= "11111111";  -- 12D5 = FF
      when "1001011010110" =>  data <= "11111111";  -- 12D6 = FF
      when "1001011010111" =>  data <= "11111111";  -- 12D7 = FF
      when "1001011011000" =>  data <= "11111111";  -- 12D8 = FF
      when "1001011011001" =>  data <= "11111111";  -- 12D9 = FF
      when "1001011011010" =>  data <= "11111111";  -- 12DA = FF
      when "1001011011011" =>  data <= "11111111";  -- 12DB = FF
      when "1001011011100" =>  data <= "11111111";  -- 12DC = FF
      when "1001011011101" =>  data <= "11111111";  -- 12DD = FF
      when "1001011011110" =>  data <= "11111111";  -- 12DE = FF
      when "1001011011111" =>  data <= "11111111";  -- 12DF = FF
      when "1001011100000" =>  data <= "11111111";  -- 12E0 = FF
      when "1001011100001" =>  data <= "11111111";  -- 12E1 = FF
      when "1001011100010" =>  data <= "11111111";  -- 12E2 = FF
      when "1001011100011" =>  data <= "11111111";  -- 12E3 = FF
      when "1001011100100" =>  data <= "11111111";  -- 12E4 = FF
      when "1001011100101" =>  data <= "11111111";  -- 12E5 = FF
      when "1001011100110" =>  data <= "11111111";  -- 12E6 = FF
      when "1001011100111" =>  data <= "11111111";  -- 12E7 = FF
      when "1001011101000" =>  data <= "11111111";  -- 12E8 = FF
      when "1001011101001" =>  data <= "11111111";  -- 12E9 = FF
      when "1001011101010" =>  data <= "11111111";  -- 12EA = FF
      when "1001011101011" =>  data <= "11111111";  -- 12EB = FF
      when "1001011101100" =>  data <= "11111111";  -- 12EC = FF
      when "1001011101101" =>  data <= "11111111";  -- 12ED = FF
      when "1001011101110" =>  data <= "11111111";  -- 12EE = FF
      when "1001011101111" =>  data <= "11111111";  -- 12EF = FF
      when "1001011110000" =>  data <= "11111111";  -- 12F0 = FF
      when "1001011110001" =>  data <= "11111111";  -- 12F1 = FF
      when "1001011110010" =>  data <= "11111111";  -- 12F2 = FF
      when "1001011110011" =>  data <= "11111111";  -- 12F3 = FF
      when "1001011110100" =>  data <= "11111111";  -- 12F4 = FF
      when "1001011110101" =>  data <= "11111111";  -- 12F5 = FF
      when "1001011110110" =>  data <= "11111111";  -- 12F6 = FF
      when "1001011110111" =>  data <= "11111111";  -- 12F7 = FF
      when "1001011111000" =>  data <= "11111111";  -- 12F8 = FF
      when "1001011111001" =>  data <= "11111111";  -- 12F9 = FF
      when "1001011111010" =>  data <= "11111111";  -- 12FA = FF
      when "1001011111011" =>  data <= "11111111";  -- 12FB = FF
      when "1001011111100" =>  data <= "11111111";  -- 12FC = FF
      when "1001011111101" =>  data <= "11111111";  -- 12FD = FF
      when "1001011111110" =>  data <= "11111111";  -- 12FE = FF
      when "1001011111111" =>  data <= "11111111";  -- 12FF = FF
      when "1001100000000" =>  data <= "11111111";  -- 1300 = FF
      when "1001100000001" =>  data <= "11111111";  -- 1301 = FF
      when "1001100000010" =>  data <= "11111111";  -- 1302 = FF
      when "1001100000011" =>  data <= "11111111";  -- 1303 = FF
      when "1001100000100" =>  data <= "11111111";  -- 1304 = FF
      when "1001100000101" =>  data <= "11111111";  -- 1305 = FF
      when "1001100000110" =>  data <= "11111111";  -- 1306 = FF
      when "1001100000111" =>  data <= "11111111";  -- 1307 = FF
      when "1001100001000" =>  data <= "11111111";  -- 1308 = FF
      when "1001100001001" =>  data <= "11111111";  -- 1309 = FF
      when "1001100001010" =>  data <= "11111111";  -- 130A = FF
      when "1001100001011" =>  data <= "11111111";  -- 130B = FF
      when "1001100001100" =>  data <= "11111111";  -- 130C = FF
      when "1001100001101" =>  data <= "11111111";  -- 130D = FF
      when "1001100001110" =>  data <= "11111111";  -- 130E = FF
      when "1001100001111" =>  data <= "11111111";  -- 130F = FF
      when "1001100010000" =>  data <= "11111111";  -- 1310 = FF
      when "1001100010001" =>  data <= "11111111";  -- 1311 = FF
      when "1001100010010" =>  data <= "11111111";  -- 1312 = FF
      when "1001100010011" =>  data <= "11111111";  -- 1313 = FF
      when "1001100010100" =>  data <= "11111111";  -- 1314 = FF
      when "1001100010101" =>  data <= "11111111";  -- 1315 = FF
      when "1001100010110" =>  data <= "11111111";  -- 1316 = FF
      when "1001100010111" =>  data <= "11111111";  -- 1317 = FF
      when "1001100011000" =>  data <= "11111111";  -- 1318 = FF
      when "1001100011001" =>  data <= "11111111";  -- 1319 = FF
      when "1001100011010" =>  data <= "11111111";  -- 131A = FF
      when "1001100011011" =>  data <= "11111111";  -- 131B = FF
      when "1001100011100" =>  data <= "11111111";  -- 131C = FF
      when "1001100011101" =>  data <= "11111111";  -- 131D = FF
      when "1001100011110" =>  data <= "11111111";  -- 131E = FF
      when "1001100011111" =>  data <= "11111111";  -- 131F = FF
      when "1001100100000" =>  data <= "11111111";  -- 1320 = FF
      when "1001100100001" =>  data <= "11111111";  -- 1321 = FF
      when "1001100100010" =>  data <= "11111111";  -- 1322 = FF
      when "1001100100011" =>  data <= "11111111";  -- 1323 = FF
      when "1001100100100" =>  data <= "11111111";  -- 1324 = FF
      when "1001100100101" =>  data <= "11111111";  -- 1325 = FF
      when "1001100100110" =>  data <= "11111111";  -- 1326 = FF
      when "1001100100111" =>  data <= "11111111";  -- 1327 = FF
      when "1001100101000" =>  data <= "11111111";  -- 1328 = FF
      when "1001100101001" =>  data <= "11111111";  -- 1329 = FF
      when "1001100101010" =>  data <= "11111111";  -- 132A = FF
      when "1001100101011" =>  data <= "11111111";  -- 132B = FF
      when "1001100101100" =>  data <= "11111111";  -- 132C = FF
      when "1001100101101" =>  data <= "11111111";  -- 132D = FF
      when "1001100101110" =>  data <= "11111111";  -- 132E = FF
      when "1001100101111" =>  data <= "11111111";  -- 132F = FF
      when "1001100110000" =>  data <= "11111111";  -- 1330 = FF
      when "1001100110001" =>  data <= "11111111";  -- 1331 = FF
      when "1001100110010" =>  data <= "11111111";  -- 1332 = FF
      when "1001100110011" =>  data <= "11111111";  -- 1333 = FF
      when "1001100110100" =>  data <= "11111111";  -- 1334 = FF
      when "1001100110101" =>  data <= "11111111";  -- 1335 = FF
      when "1001100110110" =>  data <= "11111111";  -- 1336 = FF
      when "1001100110111" =>  data <= "11111111";  -- 1337 = FF
      when "1001100111000" =>  data <= "11111111";  -- 1338 = FF
      when "1001100111001" =>  data <= "11111111";  -- 1339 = FF
      when "1001100111010" =>  data <= "11111111";  -- 133A = FF
      when "1001100111011" =>  data <= "11111111";  -- 133B = FF
      when "1001100111100" =>  data <= "11111111";  -- 133C = FF
      when "1001100111101" =>  data <= "11111111";  -- 133D = FF
      when "1001100111110" =>  data <= "11111111";  -- 133E = FF
      when "1001100111111" =>  data <= "11111111";  -- 133F = FF
      when "1001101000000" =>  data <= "11111111";  -- 1340 = FF
      when "1001101000001" =>  data <= "11111111";  -- 1341 = FF
      when "1001101000010" =>  data <= "11111111";  -- 1342 = FF
      when "1001101000011" =>  data <= "11111111";  -- 1343 = FF
      when "1001101000100" =>  data <= "11111111";  -- 1344 = FF
      when "1001101000101" =>  data <= "11111111";  -- 1345 = FF
      when "1001101000110" =>  data <= "11111111";  -- 1346 = FF
      when "1001101000111" =>  data <= "11111111";  -- 1347 = FF
      when "1001101001000" =>  data <= "11111111";  -- 1348 = FF
      when "1001101001001" =>  data <= "11111111";  -- 1349 = FF
      when "1001101001010" =>  data <= "11111111";  -- 134A = FF
      when "1001101001011" =>  data <= "11111111";  -- 134B = FF
      when "1001101001100" =>  data <= "11111111";  -- 134C = FF
      when "1001101001101" =>  data <= "11111111";  -- 134D = FF
      when "1001101001110" =>  data <= "11111111";  -- 134E = FF
      when "1001101001111" =>  data <= "11111111";  -- 134F = FF
      when "1001101010000" =>  data <= "11111111";  -- 1350 = FF
      when "1001101010001" =>  data <= "11111111";  -- 1351 = FF
      when "1001101010010" =>  data <= "11111111";  -- 1352 = FF
      when "1001101010011" =>  data <= "11111111";  -- 1353 = FF
      when "1001101010100" =>  data <= "11111111";  -- 1354 = FF
      when "1001101010101" =>  data <= "11111111";  -- 1355 = FF
      when "1001101010110" =>  data <= "11111111";  -- 1356 = FF
      when "1001101010111" =>  data <= "11111111";  -- 1357 = FF
      when "1001101011000" =>  data <= "11111111";  -- 1358 = FF
      when "1001101011001" =>  data <= "11111111";  -- 1359 = FF
      when "1001101011010" =>  data <= "11111111";  -- 135A = FF
      when "1001101011011" =>  data <= "11111111";  -- 135B = FF
      when "1001101011100" =>  data <= "11111111";  -- 135C = FF
      when "1001101011101" =>  data <= "11111111";  -- 135D = FF
      when "1001101011110" =>  data <= "11111111";  -- 135E = FF
      when "1001101011111" =>  data <= "11111111";  -- 135F = FF
      when "1001101100000" =>  data <= "11111111";  -- 1360 = FF
      when "1001101100001" =>  data <= "11111111";  -- 1361 = FF
      when "1001101100010" =>  data <= "11111111";  -- 1362 = FF
      when "1001101100011" =>  data <= "11111111";  -- 1363 = FF
      when "1001101100100" =>  data <= "11111111";  -- 1364 = FF
      when "1001101100101" =>  data <= "11111111";  -- 1365 = FF
      when "1001101100110" =>  data <= "11111111";  -- 1366 = FF
      when "1001101100111" =>  data <= "11111111";  -- 1367 = FF
      when "1001101101000" =>  data <= "11111111";  -- 1368 = FF
      when "1001101101001" =>  data <= "11111111";  -- 1369 = FF
      when "1001101101010" =>  data <= "11111111";  -- 136A = FF
      when "1001101101011" =>  data <= "11111111";  -- 136B = FF
      when "1001101101100" =>  data <= "11111111";  -- 136C = FF
      when "1001101101101" =>  data <= "11111111";  -- 136D = FF
      when "1001101101110" =>  data <= "11111111";  -- 136E = FF
      when "1001101101111" =>  data <= "11111111";  -- 136F = FF
      when "1001101110000" =>  data <= "11111111";  -- 1370 = FF
      when "1001101110001" =>  data <= "11111111";  -- 1371 = FF
      when "1001101110010" =>  data <= "11111111";  -- 1372 = FF
      when "1001101110011" =>  data <= "11111111";  -- 1373 = FF
      when "1001101110100" =>  data <= "11111111";  -- 1374 = FF
      when "1001101110101" =>  data <= "11111111";  -- 1375 = FF
      when "1001101110110" =>  data <= "11111111";  -- 1376 = FF
      when "1001101110111" =>  data <= "11111111";  -- 1377 = FF
      when "1001101111000" =>  data <= "11111111";  -- 1378 = FF
      when "1001101111001" =>  data <= "11111111";  -- 1379 = FF
      when "1001101111010" =>  data <= "11111111";  -- 137A = FF
      when "1001101111011" =>  data <= "11111111";  -- 137B = FF
      when "1001101111100" =>  data <= "11111111";  -- 137C = FF
      when "1001101111101" =>  data <= "11111111";  -- 137D = FF
      when "1001101111110" =>  data <= "11111111";  -- 137E = FF
      when "1001101111111" =>  data <= "11111111";  -- 137F = FF
      when "1001110000000" =>  data <= "11111111";  -- 1380 = FF
      when "1001110000001" =>  data <= "11111111";  -- 1381 = FF
      when "1001110000010" =>  data <= "11111111";  -- 1382 = FF
      when "1001110000011" =>  data <= "11111111";  -- 1383 = FF
      when "1001110000100" =>  data <= "11111111";  -- 1384 = FF
      when "1001110000101" =>  data <= "11111111";  -- 1385 = FF
      when "1001110000110" =>  data <= "11111111";  -- 1386 = FF
      when "1001110000111" =>  data <= "11111111";  -- 1387 = FF
      when "1001110001000" =>  data <= "11111111";  -- 1388 = FF
      when "1001110001001" =>  data <= "11111111";  -- 1389 = FF
      when "1001110001010" =>  data <= "11111111";  -- 138A = FF
      when "1001110001011" =>  data <= "11111111";  -- 138B = FF
      when "1001110001100" =>  data <= "11111111";  -- 138C = FF
      when "1001110001101" =>  data <= "11111111";  -- 138D = FF
      when "1001110001110" =>  data <= "11111111";  -- 138E = FF
      when "1001110001111" =>  data <= "11111111";  -- 138F = FF
      when "1001110010000" =>  data <= "11111111";  -- 1390 = FF
      when "1001110010001" =>  data <= "11111111";  -- 1391 = FF
      when "1001110010010" =>  data <= "11111111";  -- 1392 = FF
      when "1001110010011" =>  data <= "11111111";  -- 1393 = FF
      when "1001110010100" =>  data <= "11111111";  -- 1394 = FF
      when "1001110010101" =>  data <= "11111111";  -- 1395 = FF
      when "1001110010110" =>  data <= "11111111";  -- 1396 = FF
      when "1001110010111" =>  data <= "11111111";  -- 1397 = FF
      when "1001110011000" =>  data <= "11111111";  -- 1398 = FF
      when "1001110011001" =>  data <= "11111111";  -- 1399 = FF
      when "1001110011010" =>  data <= "11111111";  -- 139A = FF
      when "1001110011011" =>  data <= "11111111";  -- 139B = FF
      when "1001110011100" =>  data <= "11111111";  -- 139C = FF
      when "1001110011101" =>  data <= "11111111";  -- 139D = FF
      when "1001110011110" =>  data <= "11111111";  -- 139E = FF
      when "1001110011111" =>  data <= "11111111";  -- 139F = FF
      when "1001110100000" =>  data <= "11111111";  -- 13A0 = FF
      when "1001110100001" =>  data <= "11111111";  -- 13A1 = FF
      when "1001110100010" =>  data <= "11111111";  -- 13A2 = FF
      when "1001110100011" =>  data <= "11111111";  -- 13A3 = FF
      when "1001110100100" =>  data <= "11111111";  -- 13A4 = FF
      when "1001110100101" =>  data <= "11111111";  -- 13A5 = FF
      when "1001110100110" =>  data <= "11111111";  -- 13A6 = FF
      when "1001110100111" =>  data <= "11111111";  -- 13A7 = FF
      when "1001110101000" =>  data <= "11111111";  -- 13A8 = FF
      when "1001110101001" =>  data <= "11111111";  -- 13A9 = FF
      when "1001110101010" =>  data <= "11111111";  -- 13AA = FF
      when "1001110101011" =>  data <= "11111111";  -- 13AB = FF
      when "1001110101100" =>  data <= "11111111";  -- 13AC = FF
      when "1001110101101" =>  data <= "11111111";  -- 13AD = FF
      when "1001110101110" =>  data <= "11111111";  -- 13AE = FF
      when "1001110101111" =>  data <= "11111111";  -- 13AF = FF
      when "1001110110000" =>  data <= "11111111";  -- 13B0 = FF
      when "1001110110001" =>  data <= "11111111";  -- 13B1 = FF
      when "1001110110010" =>  data <= "11111111";  -- 13B2 = FF
      when "1001110110011" =>  data <= "11111111";  -- 13B3 = FF
      when "1001110110100" =>  data <= "11111111";  -- 13B4 = FF
      when "1001110110101" =>  data <= "11111111";  -- 13B5 = FF
      when "1001110110110" =>  data <= "11111111";  -- 13B6 = FF
      when "1001110110111" =>  data <= "11111111";  -- 13B7 = FF
      when "1001110111000" =>  data <= "11111111";  -- 13B8 = FF
      when "1001110111001" =>  data <= "11111111";  -- 13B9 = FF
      when "1001110111010" =>  data <= "11111111";  -- 13BA = FF
      when "1001110111011" =>  data <= "11111111";  -- 13BB = FF
      when "1001110111100" =>  data <= "11111111";  -- 13BC = FF
      when "1001110111101" =>  data <= "11111111";  -- 13BD = FF
      when "1001110111110" =>  data <= "11111111";  -- 13BE = FF
      when "1001110111111" =>  data <= "11111111";  -- 13BF = FF
      when "1001111000000" =>  data <= "11111111";  -- 13C0 = FF
      when "1001111000001" =>  data <= "11111111";  -- 13C1 = FF
      when "1001111000010" =>  data <= "11111111";  -- 13C2 = FF
      when "1001111000011" =>  data <= "11111111";  -- 13C3 = FF
      when "1001111000100" =>  data <= "11111111";  -- 13C4 = FF
      when "1001111000101" =>  data <= "11111111";  -- 13C5 = FF
      when "1001111000110" =>  data <= "11111111";  -- 13C6 = FF
      when "1001111000111" =>  data <= "11111111";  -- 13C7 = FF
      when "1001111001000" =>  data <= "11111111";  -- 13C8 = FF
      when "1001111001001" =>  data <= "11111111";  -- 13C9 = FF
      when "1001111001010" =>  data <= "11111111";  -- 13CA = FF
      when "1001111001011" =>  data <= "11111111";  -- 13CB = FF
      when "1001111001100" =>  data <= "11111111";  -- 13CC = FF
      when "1001111001101" =>  data <= "11111111";  -- 13CD = FF
      when "1001111001110" =>  data <= "11111111";  -- 13CE = FF
      when "1001111001111" =>  data <= "11111111";  -- 13CF = FF
      when "1001111010000" =>  data <= "11111111";  -- 13D0 = FF
      when "1001111010001" =>  data <= "11111111";  -- 13D1 = FF
      when "1001111010010" =>  data <= "11111111";  -- 13D2 = FF
      when "1001111010011" =>  data <= "11111111";  -- 13D3 = FF
      when "1001111010100" =>  data <= "11111111";  -- 13D4 = FF
      when "1001111010101" =>  data <= "11111111";  -- 13D5 = FF
      when "1001111010110" =>  data <= "11111111";  -- 13D6 = FF
      when "1001111010111" =>  data <= "11111111";  -- 13D7 = FF
      when "1001111011000" =>  data <= "11111111";  -- 13D8 = FF
      when "1001111011001" =>  data <= "11111111";  -- 13D9 = FF
      when "1001111011010" =>  data <= "11111111";  -- 13DA = FF
      when "1001111011011" =>  data <= "11111111";  -- 13DB = FF
      when "1001111011100" =>  data <= "11111111";  -- 13DC = FF
      when "1001111011101" =>  data <= "11111111";  -- 13DD = FF
      when "1001111011110" =>  data <= "11111111";  -- 13DE = FF
      when "1001111011111" =>  data <= "11111111";  -- 13DF = FF
      when "1001111100000" =>  data <= "11111111";  -- 13E0 = FF
      when "1001111100001" =>  data <= "11111111";  -- 13E1 = FF
      when "1001111100010" =>  data <= "11111111";  -- 13E2 = FF
      when "1001111100011" =>  data <= "11111111";  -- 13E3 = FF
      when "1001111100100" =>  data <= "11111111";  -- 13E4 = FF
      when "1001111100101" =>  data <= "11111111";  -- 13E5 = FF
      when "1001111100110" =>  data <= "11111111";  -- 13E6 = FF
      when "1001111100111" =>  data <= "11111111";  -- 13E7 = FF
      when "1001111101000" =>  data <= "11111111";  -- 13E8 = FF
      when "1001111101001" =>  data <= "11111111";  -- 13E9 = FF
      when "1001111101010" =>  data <= "11111111";  -- 13EA = FF
      when "1001111101011" =>  data <= "11111111";  -- 13EB = FF
      when "1001111101100" =>  data <= "11111111";  -- 13EC = FF
      when "1001111101101" =>  data <= "11111111";  -- 13ED = FF
      when "1001111101110" =>  data <= "11111111";  -- 13EE = FF
      when "1001111101111" =>  data <= "11111111";  -- 13EF = FF
      when "1001111110000" =>  data <= "11111111";  -- 13F0 = FF
      when "1001111110001" =>  data <= "11111111";  -- 13F1 = FF
      when "1001111110010" =>  data <= "11111111";  -- 13F2 = FF
      when "1001111110011" =>  data <= "11111111";  -- 13F3 = FF
      when "1001111110100" =>  data <= "11111111";  -- 13F4 = FF
      when "1001111110101" =>  data <= "11111111";  -- 13F5 = FF
      when "1001111110110" =>  data <= "11111111";  -- 13F6 = FF
      when "1001111110111" =>  data <= "11111111";  -- 13F7 = FF
      when "1001111111000" =>  data <= "11111111";  -- 13F8 = FF
      when "1001111111001" =>  data <= "11111111";  -- 13F9 = FF
      when "1001111111010" =>  data <= "11111111";  -- 13FA = FF
      when "1001111111011" =>  data <= "11111111";  -- 13FB = FF
      when "1001111111100" =>  data <= "11111111";  -- 13FC = FF
      when "1001111111101" =>  data <= "11111111";  -- 13FD = FF
      when "1001111111110" =>  data <= "11111111";  -- 13FE = FF
      when "1001111111111" =>  data <= "11111111";  -- 13FF = FF
      when "1010000000000" =>  data <= "11111111";  -- 1400 = FF
      when "1010000000001" =>  data <= "11111111";  -- 1401 = FF
      when "1010000000010" =>  data <= "11111111";  -- 1402 = FF
      when "1010000000011" =>  data <= "11111111";  -- 1403 = FF
      when "1010000000100" =>  data <= "11111111";  -- 1404 = FF
      when "1010000000101" =>  data <= "11111111";  -- 1405 = FF
      when "1010000000110" =>  data <= "11111111";  -- 1406 = FF
      when "1010000000111" =>  data <= "11111111";  -- 1407 = FF
      when "1010000001000" =>  data <= "11111111";  -- 1408 = FF
      when "1010000001001" =>  data <= "11111111";  -- 1409 = FF
      when "1010000001010" =>  data <= "11111111";  -- 140A = FF
      when "1010000001011" =>  data <= "11111111";  -- 140B = FF
      when "1010000001100" =>  data <= "11111111";  -- 140C = FF
      when "1010000001101" =>  data <= "11111111";  -- 140D = FF
      when "1010000001110" =>  data <= "11111111";  -- 140E = FF
      when "1010000001111" =>  data <= "11111111";  -- 140F = FF
      when "1010000010000" =>  data <= "11111111";  -- 1410 = FF
      when "1010000010001" =>  data <= "11111111";  -- 1411 = FF
      when "1010000010010" =>  data <= "11111111";  -- 1412 = FF
      when "1010000010011" =>  data <= "11111111";  -- 1413 = FF
      when "1010000010100" =>  data <= "11111111";  -- 1414 = FF
      when "1010000010101" =>  data <= "11111111";  -- 1415 = FF
      when "1010000010110" =>  data <= "11111111";  -- 1416 = FF
      when "1010000010111" =>  data <= "11111111";  -- 1417 = FF
      when "1010000011000" =>  data <= "11111111";  -- 1418 = FF
      when "1010000011001" =>  data <= "11111111";  -- 1419 = FF
      when "1010000011010" =>  data <= "11111111";  -- 141A = FF
      when "1010000011011" =>  data <= "11111111";  -- 141B = FF
      when "1010000011100" =>  data <= "11111111";  -- 141C = FF
      when "1010000011101" =>  data <= "11111111";  -- 141D = FF
      when "1010000011110" =>  data <= "11111111";  -- 141E = FF
      when "1010000011111" =>  data <= "11111111";  -- 141F = FF
      when "1010000100000" =>  data <= "11111111";  -- 1420 = FF
      when "1010000100001" =>  data <= "11111111";  -- 1421 = FF
      when "1010000100010" =>  data <= "11111111";  -- 1422 = FF
      when "1010000100011" =>  data <= "11111111";  -- 1423 = FF
      when "1010000100100" =>  data <= "11111111";  -- 1424 = FF
      when "1010000100101" =>  data <= "11111111";  -- 1425 = FF
      when "1010000100110" =>  data <= "11111111";  -- 1426 = FF
      when "1010000100111" =>  data <= "11111111";  -- 1427 = FF
      when "1010000101000" =>  data <= "11111111";  -- 1428 = FF
      when "1010000101001" =>  data <= "11111111";  -- 1429 = FF
      when "1010000101010" =>  data <= "11111111";  -- 142A = FF
      when "1010000101011" =>  data <= "11111111";  -- 142B = FF
      when "1010000101100" =>  data <= "11111111";  -- 142C = FF
      when "1010000101101" =>  data <= "11111111";  -- 142D = FF
      when "1010000101110" =>  data <= "11111111";  -- 142E = FF
      when "1010000101111" =>  data <= "11111111";  -- 142F = FF
      when "1010000110000" =>  data <= "11111111";  -- 1430 = FF
      when "1010000110001" =>  data <= "11111111";  -- 1431 = FF
      when "1010000110010" =>  data <= "11111111";  -- 1432 = FF
      when "1010000110011" =>  data <= "11111111";  -- 1433 = FF
      when "1010000110100" =>  data <= "11111111";  -- 1434 = FF
      when "1010000110101" =>  data <= "11111111";  -- 1435 = FF
      when "1010000110110" =>  data <= "11111111";  -- 1436 = FF
      when "1010000110111" =>  data <= "11111111";  -- 1437 = FF
      when "1010000111000" =>  data <= "11111111";  -- 1438 = FF
      when "1010000111001" =>  data <= "11111111";  -- 1439 = FF
      when "1010000111010" =>  data <= "11111111";  -- 143A = FF
      when "1010000111011" =>  data <= "11111111";  -- 143B = FF
      when "1010000111100" =>  data <= "11111111";  -- 143C = FF
      when "1010000111101" =>  data <= "11111111";  -- 143D = FF
      when "1010000111110" =>  data <= "11111111";  -- 143E = FF
      when "1010000111111" =>  data <= "11111111";  -- 143F = FF
      when "1010001000000" =>  data <= "11111111";  -- 1440 = FF
      when "1010001000001" =>  data <= "11111111";  -- 1441 = FF
      when "1010001000010" =>  data <= "11111111";  -- 1442 = FF
      when "1010001000011" =>  data <= "11111111";  -- 1443 = FF
      when "1010001000100" =>  data <= "11111111";  -- 1444 = FF
      when "1010001000101" =>  data <= "11111111";  -- 1445 = FF
      when "1010001000110" =>  data <= "11111111";  -- 1446 = FF
      when "1010001000111" =>  data <= "11111111";  -- 1447 = FF
      when "1010001001000" =>  data <= "11111111";  -- 1448 = FF
      when "1010001001001" =>  data <= "11111111";  -- 1449 = FF
      when "1010001001010" =>  data <= "11111111";  -- 144A = FF
      when "1010001001011" =>  data <= "11111111";  -- 144B = FF
      when "1010001001100" =>  data <= "11111111";  -- 144C = FF
      when "1010001001101" =>  data <= "11111111";  -- 144D = FF
      when "1010001001110" =>  data <= "11111111";  -- 144E = FF
      when "1010001001111" =>  data <= "11111111";  -- 144F = FF
      when "1010001010000" =>  data <= "11111111";  -- 1450 = FF
      when "1010001010001" =>  data <= "11111111";  -- 1451 = FF
      when "1010001010010" =>  data <= "11111111";  -- 1452 = FF
      when "1010001010011" =>  data <= "11111111";  -- 1453 = FF
      when "1010001010100" =>  data <= "11111111";  -- 1454 = FF
      when "1010001010101" =>  data <= "11111111";  -- 1455 = FF
      when "1010001010110" =>  data <= "11111111";  -- 1456 = FF
      when "1010001010111" =>  data <= "11111111";  -- 1457 = FF
      when "1010001011000" =>  data <= "11111111";  -- 1458 = FF
      when "1010001011001" =>  data <= "11111111";  -- 1459 = FF
      when "1010001011010" =>  data <= "11111111";  -- 145A = FF
      when "1010001011011" =>  data <= "11111111";  -- 145B = FF
      when "1010001011100" =>  data <= "11111111";  -- 145C = FF
      when "1010001011101" =>  data <= "11111111";  -- 145D = FF
      when "1010001011110" =>  data <= "11111111";  -- 145E = FF
      when "1010001011111" =>  data <= "11111111";  -- 145F = FF
      when "1010001100000" =>  data <= "11111111";  -- 1460 = FF
      when "1010001100001" =>  data <= "11111111";  -- 1461 = FF
      when "1010001100010" =>  data <= "11111111";  -- 1462 = FF
      when "1010001100011" =>  data <= "11111111";  -- 1463 = FF
      when "1010001100100" =>  data <= "11111111";  -- 1464 = FF
      when "1010001100101" =>  data <= "11111111";  -- 1465 = FF
      when "1010001100110" =>  data <= "11111111";  -- 1466 = FF
      when "1010001100111" =>  data <= "11111111";  -- 1467 = FF
      when "1010001101000" =>  data <= "11111111";  -- 1468 = FF
      when "1010001101001" =>  data <= "11111111";  -- 1469 = FF
      when "1010001101010" =>  data <= "11111111";  -- 146A = FF
      when "1010001101011" =>  data <= "11111111";  -- 146B = FF
      when "1010001101100" =>  data <= "11111111";  -- 146C = FF
      when "1010001101101" =>  data <= "11111111";  -- 146D = FF
      when "1010001101110" =>  data <= "11111111";  -- 146E = FF
      when "1010001101111" =>  data <= "11111111";  -- 146F = FF
      when "1010001110000" =>  data <= "11111111";  -- 1470 = FF
      when "1010001110001" =>  data <= "11111111";  -- 1471 = FF
      when "1010001110010" =>  data <= "11111111";  -- 1472 = FF
      when "1010001110011" =>  data <= "11111111";  -- 1473 = FF
      when "1010001110100" =>  data <= "11111111";  -- 1474 = FF
      when "1010001110101" =>  data <= "11111111";  -- 1475 = FF
      when "1010001110110" =>  data <= "11111111";  -- 1476 = FF
      when "1010001110111" =>  data <= "11111111";  -- 1477 = FF
      when "1010001111000" =>  data <= "11111111";  -- 1478 = FF
      when "1010001111001" =>  data <= "11111111";  -- 1479 = FF
      when "1010001111010" =>  data <= "11111111";  -- 147A = FF
      when "1010001111011" =>  data <= "11111111";  -- 147B = FF
      when "1010001111100" =>  data <= "11111111";  -- 147C = FF
      when "1010001111101" =>  data <= "11111111";  -- 147D = FF
      when "1010001111110" =>  data <= "11111111";  -- 147E = FF
      when "1010001111111" =>  data <= "11111111";  -- 147F = FF
      when "1010010000000" =>  data <= "11111111";  -- 1480 = FF
      when "1010010000001" =>  data <= "11111111";  -- 1481 = FF
      when "1010010000010" =>  data <= "11111111";  -- 1482 = FF
      when "1010010000011" =>  data <= "11111111";  -- 1483 = FF
      when "1010010000100" =>  data <= "11111111";  -- 1484 = FF
      when "1010010000101" =>  data <= "11111111";  -- 1485 = FF
      when "1010010000110" =>  data <= "11111111";  -- 1486 = FF
      when "1010010000111" =>  data <= "11111111";  -- 1487 = FF
      when "1010010001000" =>  data <= "11111111";  -- 1488 = FF
      when "1010010001001" =>  data <= "11111111";  -- 1489 = FF
      when "1010010001010" =>  data <= "11111111";  -- 148A = FF
      when "1010010001011" =>  data <= "11111111";  -- 148B = FF
      when "1010010001100" =>  data <= "11111111";  -- 148C = FF
      when "1010010001101" =>  data <= "11111111";  -- 148D = FF
      when "1010010001110" =>  data <= "11111111";  -- 148E = FF
      when "1010010001111" =>  data <= "11111111";  -- 148F = FF
      when "1010010010000" =>  data <= "11111111";  -- 1490 = FF
      when "1010010010001" =>  data <= "11111111";  -- 1491 = FF
      when "1010010010010" =>  data <= "11111111";  -- 1492 = FF
      when "1010010010011" =>  data <= "11111111";  -- 1493 = FF
      when "1010010010100" =>  data <= "11111111";  -- 1494 = FF
      when "1010010010101" =>  data <= "11111111";  -- 1495 = FF
      when "1010010010110" =>  data <= "11111111";  -- 1496 = FF
      when "1010010010111" =>  data <= "11111111";  -- 1497 = FF
      when "1010010011000" =>  data <= "11111111";  -- 1498 = FF
      when "1010010011001" =>  data <= "11111111";  -- 1499 = FF
      when "1010010011010" =>  data <= "11111111";  -- 149A = FF
      when "1010010011011" =>  data <= "11111111";  -- 149B = FF
      when "1010010011100" =>  data <= "11111111";  -- 149C = FF
      when "1010010011101" =>  data <= "11111111";  -- 149D = FF
      when "1010010011110" =>  data <= "11111111";  -- 149E = FF
      when "1010010011111" =>  data <= "11111111";  -- 149F = FF
      when "1010010100000" =>  data <= "11111111";  -- 14A0 = FF
      when "1010010100001" =>  data <= "11111111";  -- 14A1 = FF
      when "1010010100010" =>  data <= "11111111";  -- 14A2 = FF
      when "1010010100011" =>  data <= "11111111";  -- 14A3 = FF
      when "1010010100100" =>  data <= "11111111";  -- 14A4 = FF
      when "1010010100101" =>  data <= "11111111";  -- 14A5 = FF
      when "1010010100110" =>  data <= "11111111";  -- 14A6 = FF
      when "1010010100111" =>  data <= "11111111";  -- 14A7 = FF
      when "1010010101000" =>  data <= "11111111";  -- 14A8 = FF
      when "1010010101001" =>  data <= "11111111";  -- 14A9 = FF
      when "1010010101010" =>  data <= "11111111";  -- 14AA = FF
      when "1010010101011" =>  data <= "11111111";  -- 14AB = FF
      when "1010010101100" =>  data <= "11111111";  -- 14AC = FF
      when "1010010101101" =>  data <= "11111111";  -- 14AD = FF
      when "1010010101110" =>  data <= "11111111";  -- 14AE = FF
      when "1010010101111" =>  data <= "11111111";  -- 14AF = FF
      when "1010010110000" =>  data <= "11111111";  -- 14B0 = FF
      when "1010010110001" =>  data <= "11111111";  -- 14B1 = FF
      when "1010010110010" =>  data <= "11111111";  -- 14B2 = FF
      when "1010010110011" =>  data <= "11111111";  -- 14B3 = FF
      when "1010010110100" =>  data <= "11111111";  -- 14B4 = FF
      when "1010010110101" =>  data <= "11111111";  -- 14B5 = FF
      when "1010010110110" =>  data <= "11111111";  -- 14B6 = FF
      when "1010010110111" =>  data <= "11111111";  -- 14B7 = FF
      when "1010010111000" =>  data <= "11111111";  -- 14B8 = FF
      when "1010010111001" =>  data <= "11111111";  -- 14B9 = FF
      when "1010010111010" =>  data <= "11111111";  -- 14BA = FF
      when "1010010111011" =>  data <= "11111111";  -- 14BB = FF
      when "1010010111100" =>  data <= "11111111";  -- 14BC = FF
      when "1010010111101" =>  data <= "11111111";  -- 14BD = FF
      when "1010010111110" =>  data <= "11111111";  -- 14BE = FF
      when "1010010111111" =>  data <= "11111111";  -- 14BF = FF
      when "1010011000000" =>  data <= "11111111";  -- 14C0 = FF
      when "1010011000001" =>  data <= "11111111";  -- 14C1 = FF
      when "1010011000010" =>  data <= "11111111";  -- 14C2 = FF
      when "1010011000011" =>  data <= "11111111";  -- 14C3 = FF
      when "1010011000100" =>  data <= "11111111";  -- 14C4 = FF
      when "1010011000101" =>  data <= "11111111";  -- 14C5 = FF
      when "1010011000110" =>  data <= "11111111";  -- 14C6 = FF
      when "1010011000111" =>  data <= "11111111";  -- 14C7 = FF
      when "1010011001000" =>  data <= "11111111";  -- 14C8 = FF
      when "1010011001001" =>  data <= "11111111";  -- 14C9 = FF
      when "1010011001010" =>  data <= "11111111";  -- 14CA = FF
      when "1010011001011" =>  data <= "11111111";  -- 14CB = FF
      when "1010011001100" =>  data <= "11111111";  -- 14CC = FF
      when "1010011001101" =>  data <= "11111111";  -- 14CD = FF
      when "1010011001110" =>  data <= "11111111";  -- 14CE = FF
      when "1010011001111" =>  data <= "11111111";  -- 14CF = FF
      when "1010011010000" =>  data <= "11111111";  -- 14D0 = FF
      when "1010011010001" =>  data <= "11111111";  -- 14D1 = FF
      when "1010011010010" =>  data <= "11111111";  -- 14D2 = FF
      when "1010011010011" =>  data <= "11111111";  -- 14D3 = FF
      when "1010011010100" =>  data <= "11111111";  -- 14D4 = FF
      when "1010011010101" =>  data <= "11111111";  -- 14D5 = FF
      when "1010011010110" =>  data <= "11111111";  -- 14D6 = FF
      when "1010011010111" =>  data <= "11111111";  -- 14D7 = FF
      when "1010011011000" =>  data <= "11111111";  -- 14D8 = FF
      when "1010011011001" =>  data <= "11111111";  -- 14D9 = FF
      when "1010011011010" =>  data <= "11111111";  -- 14DA = FF
      when "1010011011011" =>  data <= "11111111";  -- 14DB = FF
      when "1010011011100" =>  data <= "11111111";  -- 14DC = FF
      when "1010011011101" =>  data <= "11111111";  -- 14DD = FF
      when "1010011011110" =>  data <= "11111111";  -- 14DE = FF
      when "1010011011111" =>  data <= "11111111";  -- 14DF = FF
      when "1010011100000" =>  data <= "11111111";  -- 14E0 = FF
      when "1010011100001" =>  data <= "11111111";  -- 14E1 = FF
      when "1010011100010" =>  data <= "11111111";  -- 14E2 = FF
      when "1010011100011" =>  data <= "11111111";  -- 14E3 = FF
      when "1010011100100" =>  data <= "11111111";  -- 14E4 = FF
      when "1010011100101" =>  data <= "11111111";  -- 14E5 = FF
      when "1010011100110" =>  data <= "11111111";  -- 14E6 = FF
      when "1010011100111" =>  data <= "11111111";  -- 14E7 = FF
      when "1010011101000" =>  data <= "11111111";  -- 14E8 = FF
      when "1010011101001" =>  data <= "11111111";  -- 14E9 = FF
      when "1010011101010" =>  data <= "11111111";  -- 14EA = FF
      when "1010011101011" =>  data <= "11111111";  -- 14EB = FF
      when "1010011101100" =>  data <= "11111111";  -- 14EC = FF
      when "1010011101101" =>  data <= "11111111";  -- 14ED = FF
      when "1010011101110" =>  data <= "11111111";  -- 14EE = FF
      when "1010011101111" =>  data <= "11111111";  -- 14EF = FF
      when "1010011110000" =>  data <= "11111111";  -- 14F0 = FF
      when "1010011110001" =>  data <= "11111111";  -- 14F1 = FF
      when "1010011110010" =>  data <= "11111111";  -- 14F2 = FF
      when "1010011110011" =>  data <= "11111111";  -- 14F3 = FF
      when "1010011110100" =>  data <= "11111111";  -- 14F4 = FF
      when "1010011110101" =>  data <= "11111111";  -- 14F5 = FF
      when "1010011110110" =>  data <= "11111111";  -- 14F6 = FF
      when "1010011110111" =>  data <= "11111111";  -- 14F7 = FF
      when "1010011111000" =>  data <= "11111111";  -- 14F8 = FF
      when "1010011111001" =>  data <= "11111111";  -- 14F9 = FF
      when "1010011111010" =>  data <= "11111111";  -- 14FA = FF
      when "1010011111011" =>  data <= "11111111";  -- 14FB = FF
      when "1010011111100" =>  data <= "11111111";  -- 14FC = FF
      when "1010011111101" =>  data <= "11111111";  -- 14FD = FF
      when "1010011111110" =>  data <= "11111111";  -- 14FE = FF
      when "1010011111111" =>  data <= "11111111";  -- 14FF = FF
      when "1010100000000" =>  data <= "11111111";  -- 1500 = FF
      when "1010100000001" =>  data <= "11111111";  -- 1501 = FF
      when "1010100000010" =>  data <= "11111111";  -- 1502 = FF
      when "1010100000011" =>  data <= "11111111";  -- 1503 = FF
      when "1010100000100" =>  data <= "11111111";  -- 1504 = FF
      when "1010100000101" =>  data <= "11111111";  -- 1505 = FF
      when "1010100000110" =>  data <= "11111111";  -- 1506 = FF
      when "1010100000111" =>  data <= "11111111";  -- 1507 = FF
      when "1010100001000" =>  data <= "11111111";  -- 1508 = FF
      when "1010100001001" =>  data <= "11111111";  -- 1509 = FF
      when "1010100001010" =>  data <= "11111111";  -- 150A = FF
      when "1010100001011" =>  data <= "11111111";  -- 150B = FF
      when "1010100001100" =>  data <= "11111111";  -- 150C = FF
      when "1010100001101" =>  data <= "11111111";  -- 150D = FF
      when "1010100001110" =>  data <= "11111111";  -- 150E = FF
      when "1010100001111" =>  data <= "11111111";  -- 150F = FF
      when "1010100010000" =>  data <= "11111111";  -- 1510 = FF
      when "1010100010001" =>  data <= "11111111";  -- 1511 = FF
      when "1010100010010" =>  data <= "11111111";  -- 1512 = FF
      when "1010100010011" =>  data <= "11111111";  -- 1513 = FF
      when "1010100010100" =>  data <= "11111111";  -- 1514 = FF
      when "1010100010101" =>  data <= "11111111";  -- 1515 = FF
      when "1010100010110" =>  data <= "11111111";  -- 1516 = FF
      when "1010100010111" =>  data <= "11111111";  -- 1517 = FF
      when "1010100011000" =>  data <= "11111111";  -- 1518 = FF
      when "1010100011001" =>  data <= "11111111";  -- 1519 = FF
      when "1010100011010" =>  data <= "11111111";  -- 151A = FF
      when "1010100011011" =>  data <= "11111111";  -- 151B = FF
      when "1010100011100" =>  data <= "11111111";  -- 151C = FF
      when "1010100011101" =>  data <= "11111111";  -- 151D = FF
      when "1010100011110" =>  data <= "11111111";  -- 151E = FF
      when "1010100011111" =>  data <= "11111111";  -- 151F = FF
      when "1010100100000" =>  data <= "11111111";  -- 1520 = FF
      when "1010100100001" =>  data <= "11111111";  -- 1521 = FF
      when "1010100100010" =>  data <= "11111111";  -- 1522 = FF
      when "1010100100011" =>  data <= "11111111";  -- 1523 = FF
      when "1010100100100" =>  data <= "11111111";  -- 1524 = FF
      when "1010100100101" =>  data <= "11111111";  -- 1525 = FF
      when "1010100100110" =>  data <= "11111111";  -- 1526 = FF
      when "1010100100111" =>  data <= "11111111";  -- 1527 = FF
      when "1010100101000" =>  data <= "11111111";  -- 1528 = FF
      when "1010100101001" =>  data <= "11111111";  -- 1529 = FF
      when "1010100101010" =>  data <= "11111111";  -- 152A = FF
      when "1010100101011" =>  data <= "11111111";  -- 152B = FF
      when "1010100101100" =>  data <= "11111111";  -- 152C = FF
      when "1010100101101" =>  data <= "11111111";  -- 152D = FF
      when "1010100101110" =>  data <= "11111111";  -- 152E = FF
      when "1010100101111" =>  data <= "11111111";  -- 152F = FF
      when "1010100110000" =>  data <= "11111111";  -- 1530 = FF
      when "1010100110001" =>  data <= "11111111";  -- 1531 = FF
      when "1010100110010" =>  data <= "11111111";  -- 1532 = FF
      when "1010100110011" =>  data <= "11111111";  -- 1533 = FF
      when "1010100110100" =>  data <= "11111111";  -- 1534 = FF
      when "1010100110101" =>  data <= "11111111";  -- 1535 = FF
      when "1010100110110" =>  data <= "11111111";  -- 1536 = FF
      when "1010100110111" =>  data <= "11111111";  -- 1537 = FF
      when "1010100111000" =>  data <= "11111111";  -- 1538 = FF
      when "1010100111001" =>  data <= "11111111";  -- 1539 = FF
      when "1010100111010" =>  data <= "11111111";  -- 153A = FF
      when "1010100111011" =>  data <= "11111111";  -- 153B = FF
      when "1010100111100" =>  data <= "11111111";  -- 153C = FF
      when "1010100111101" =>  data <= "11111111";  -- 153D = FF
      when "1010100111110" =>  data <= "11111111";  -- 153E = FF
      when "1010100111111" =>  data <= "11111111";  -- 153F = FF
      when "1010101000000" =>  data <= "11111111";  -- 1540 = FF
      when "1010101000001" =>  data <= "11111111";  -- 1541 = FF
      when "1010101000010" =>  data <= "11111111";  -- 1542 = FF
      when "1010101000011" =>  data <= "11111111";  -- 1543 = FF
      when "1010101000100" =>  data <= "11111111";  -- 1544 = FF
      when "1010101000101" =>  data <= "11111111";  -- 1545 = FF
      when "1010101000110" =>  data <= "11111111";  -- 1546 = FF
      when "1010101000111" =>  data <= "11111111";  -- 1547 = FF
      when "1010101001000" =>  data <= "11111111";  -- 1548 = FF
      when "1010101001001" =>  data <= "11111111";  -- 1549 = FF
      when "1010101001010" =>  data <= "11111111";  -- 154A = FF
      when "1010101001011" =>  data <= "11111111";  -- 154B = FF
      when "1010101001100" =>  data <= "11111111";  -- 154C = FF
      when "1010101001101" =>  data <= "11111111";  -- 154D = FF
      when "1010101001110" =>  data <= "11111111";  -- 154E = FF
      when "1010101001111" =>  data <= "11111111";  -- 154F = FF
      when "1010101010000" =>  data <= "11111111";  -- 1550 = FF
      when "1010101010001" =>  data <= "11111111";  -- 1551 = FF
      when "1010101010010" =>  data <= "11111111";  -- 1552 = FF
      when "1010101010011" =>  data <= "11111111";  -- 1553 = FF
      when "1010101010100" =>  data <= "11111111";  -- 1554 = FF
      when "1010101010101" =>  data <= "11111111";  -- 1555 = FF
      when "1010101010110" =>  data <= "11111111";  -- 1556 = FF
      when "1010101010111" =>  data <= "11111111";  -- 1557 = FF
      when "1010101011000" =>  data <= "11111111";  -- 1558 = FF
      when "1010101011001" =>  data <= "11111111";  -- 1559 = FF
      when "1010101011010" =>  data <= "11111111";  -- 155A = FF
      when "1010101011011" =>  data <= "11111111";  -- 155B = FF
      when "1010101011100" =>  data <= "11111111";  -- 155C = FF
      when "1010101011101" =>  data <= "11111111";  -- 155D = FF
      when "1010101011110" =>  data <= "11111111";  -- 155E = FF
      when "1010101011111" =>  data <= "11111111";  -- 155F = FF
      when "1010101100000" =>  data <= "11111111";  -- 1560 = FF
      when "1010101100001" =>  data <= "11111111";  -- 1561 = FF
      when "1010101100010" =>  data <= "11111111";  -- 1562 = FF
      when "1010101100011" =>  data <= "11111111";  -- 1563 = FF
      when "1010101100100" =>  data <= "11111111";  -- 1564 = FF
      when "1010101100101" =>  data <= "11111111";  -- 1565 = FF
      when "1010101100110" =>  data <= "11111111";  -- 1566 = FF
      when "1010101100111" =>  data <= "11111111";  -- 1567 = FF
      when "1010101101000" =>  data <= "11111111";  -- 1568 = FF
      when "1010101101001" =>  data <= "11111111";  -- 1569 = FF
      when "1010101101010" =>  data <= "11111111";  -- 156A = FF
      when "1010101101011" =>  data <= "11111111";  -- 156B = FF
      when "1010101101100" =>  data <= "11111111";  -- 156C = FF
      when "1010101101101" =>  data <= "11111111";  -- 156D = FF
      when "1010101101110" =>  data <= "11111111";  -- 156E = FF
      when "1010101101111" =>  data <= "11111111";  -- 156F = FF
      when "1010101110000" =>  data <= "11111111";  -- 1570 = FF
      when "1010101110001" =>  data <= "11111111";  -- 1571 = FF
      when "1010101110010" =>  data <= "11111111";  -- 1572 = FF
      when "1010101110011" =>  data <= "11111111";  -- 1573 = FF
      when "1010101110100" =>  data <= "11111111";  -- 1574 = FF
      when "1010101110101" =>  data <= "11111111";  -- 1575 = FF
      when "1010101110110" =>  data <= "11111111";  -- 1576 = FF
      when "1010101110111" =>  data <= "11111111";  -- 1577 = FF
      when "1010101111000" =>  data <= "11111111";  -- 1578 = FF
      when "1010101111001" =>  data <= "11111111";  -- 1579 = FF
      when "1010101111010" =>  data <= "11111111";  -- 157A = FF
      when "1010101111011" =>  data <= "11111111";  -- 157B = FF
      when "1010101111100" =>  data <= "11111111";  -- 157C = FF
      when "1010101111101" =>  data <= "11111111";  -- 157D = FF
      when "1010101111110" =>  data <= "11111111";  -- 157E = FF
      when "1010101111111" =>  data <= "11111111";  -- 157F = FF
      when "1010110000000" =>  data <= "11111111";  -- 1580 = FF
      when "1010110000001" =>  data <= "11111111";  -- 1581 = FF
      when "1010110000010" =>  data <= "11111111";  -- 1582 = FF
      when "1010110000011" =>  data <= "11111111";  -- 1583 = FF
      when "1010110000100" =>  data <= "11111111";  -- 1584 = FF
      when "1010110000101" =>  data <= "11111111";  -- 1585 = FF
      when "1010110000110" =>  data <= "11111111";  -- 1586 = FF
      when "1010110000111" =>  data <= "11111111";  -- 1587 = FF
      when "1010110001000" =>  data <= "11111111";  -- 1588 = FF
      when "1010110001001" =>  data <= "11111111";  -- 1589 = FF
      when "1010110001010" =>  data <= "11111111";  -- 158A = FF
      when "1010110001011" =>  data <= "11111111";  -- 158B = FF
      when "1010110001100" =>  data <= "11111111";  -- 158C = FF
      when "1010110001101" =>  data <= "11111111";  -- 158D = FF
      when "1010110001110" =>  data <= "11111111";  -- 158E = FF
      when "1010110001111" =>  data <= "11111111";  -- 158F = FF
      when "1010110010000" =>  data <= "11111111";  -- 1590 = FF
      when "1010110010001" =>  data <= "11111111";  -- 1591 = FF
      when "1010110010010" =>  data <= "11111111";  -- 1592 = FF
      when "1010110010011" =>  data <= "11111111";  -- 1593 = FF
      when "1010110010100" =>  data <= "11111111";  -- 1594 = FF
      when "1010110010101" =>  data <= "11111111";  -- 1595 = FF
      when "1010110010110" =>  data <= "11111111";  -- 1596 = FF
      when "1010110010111" =>  data <= "11111111";  -- 1597 = FF
      when "1010110011000" =>  data <= "11111111";  -- 1598 = FF
      when "1010110011001" =>  data <= "11111111";  -- 1599 = FF
      when "1010110011010" =>  data <= "11111111";  -- 159A = FF
      when "1010110011011" =>  data <= "11111111";  -- 159B = FF
      when "1010110011100" =>  data <= "11111111";  -- 159C = FF
      when "1010110011101" =>  data <= "11111111";  -- 159D = FF
      when "1010110011110" =>  data <= "11111111";  -- 159E = FF
      when "1010110011111" =>  data <= "11111111";  -- 159F = FF
      when "1010110100000" =>  data <= "11111111";  -- 15A0 = FF
      when "1010110100001" =>  data <= "11111111";  -- 15A1 = FF
      when "1010110100010" =>  data <= "11111111";  -- 15A2 = FF
      when "1010110100011" =>  data <= "11111111";  -- 15A3 = FF
      when "1010110100100" =>  data <= "11111111";  -- 15A4 = FF
      when "1010110100101" =>  data <= "11111111";  -- 15A5 = FF
      when "1010110100110" =>  data <= "11111111";  -- 15A6 = FF
      when "1010110100111" =>  data <= "11111111";  -- 15A7 = FF
      when "1010110101000" =>  data <= "11111111";  -- 15A8 = FF
      when "1010110101001" =>  data <= "11111111";  -- 15A9 = FF
      when "1010110101010" =>  data <= "11111111";  -- 15AA = FF
      when "1010110101011" =>  data <= "11111111";  -- 15AB = FF
      when "1010110101100" =>  data <= "11111111";  -- 15AC = FF
      when "1010110101101" =>  data <= "11111111";  -- 15AD = FF
      when "1010110101110" =>  data <= "11111111";  -- 15AE = FF
      when "1010110101111" =>  data <= "11111111";  -- 15AF = FF
      when "1010110110000" =>  data <= "11111111";  -- 15B0 = FF
      when "1010110110001" =>  data <= "11111111";  -- 15B1 = FF
      when "1010110110010" =>  data <= "11111111";  -- 15B2 = FF
      when "1010110110011" =>  data <= "11111111";  -- 15B3 = FF
      when "1010110110100" =>  data <= "11111111";  -- 15B4 = FF
      when "1010110110101" =>  data <= "11111111";  -- 15B5 = FF
      when "1010110110110" =>  data <= "11111111";  -- 15B6 = FF
      when "1010110110111" =>  data <= "11111111";  -- 15B7 = FF
      when "1010110111000" =>  data <= "11111111";  -- 15B8 = FF
      when "1010110111001" =>  data <= "11111111";  -- 15B9 = FF
      when "1010110111010" =>  data <= "11111111";  -- 15BA = FF
      when "1010110111011" =>  data <= "11111111";  -- 15BB = FF
      when "1010110111100" =>  data <= "11111111";  -- 15BC = FF
      when "1010110111101" =>  data <= "11111111";  -- 15BD = FF
      when "1010110111110" =>  data <= "11111111";  -- 15BE = FF
      when "1010110111111" =>  data <= "11111111";  -- 15BF = FF
      when "1010111000000" =>  data <= "11111111";  -- 15C0 = FF
      when "1010111000001" =>  data <= "11111111";  -- 15C1 = FF
      when "1010111000010" =>  data <= "11111111";  -- 15C2 = FF
      when "1010111000011" =>  data <= "11111111";  -- 15C3 = FF
      when "1010111000100" =>  data <= "11111111";  -- 15C4 = FF
      when "1010111000101" =>  data <= "11111111";  -- 15C5 = FF
      when "1010111000110" =>  data <= "11111111";  -- 15C6 = FF
      when "1010111000111" =>  data <= "11111111";  -- 15C7 = FF
      when "1010111001000" =>  data <= "11111111";  -- 15C8 = FF
      when "1010111001001" =>  data <= "11111111";  -- 15C9 = FF
      when "1010111001010" =>  data <= "11111111";  -- 15CA = FF
      when "1010111001011" =>  data <= "11111111";  -- 15CB = FF
      when "1010111001100" =>  data <= "11111111";  -- 15CC = FF
      when "1010111001101" =>  data <= "11111111";  -- 15CD = FF
      when "1010111001110" =>  data <= "11111111";  -- 15CE = FF
      when "1010111001111" =>  data <= "11111111";  -- 15CF = FF
      when "1010111010000" =>  data <= "11111111";  -- 15D0 = FF
      when "1010111010001" =>  data <= "11111111";  -- 15D1 = FF
      when "1010111010010" =>  data <= "11111111";  -- 15D2 = FF
      when "1010111010011" =>  data <= "11111111";  -- 15D3 = FF
      when "1010111010100" =>  data <= "11111111";  -- 15D4 = FF
      when "1010111010101" =>  data <= "11111111";  -- 15D5 = FF
      when "1010111010110" =>  data <= "11111111";  -- 15D6 = FF
      when "1010111010111" =>  data <= "11111111";  -- 15D7 = FF
      when "1010111011000" =>  data <= "11111111";  -- 15D8 = FF
      when "1010111011001" =>  data <= "11111111";  -- 15D9 = FF
      when "1010111011010" =>  data <= "11111111";  -- 15DA = FF
      when "1010111011011" =>  data <= "11111111";  -- 15DB = FF
      when "1010111011100" =>  data <= "11111111";  -- 15DC = FF
      when "1010111011101" =>  data <= "11111111";  -- 15DD = FF
      when "1010111011110" =>  data <= "11111111";  -- 15DE = FF
      when "1010111011111" =>  data <= "11111111";  -- 15DF = FF
      when "1010111100000" =>  data <= "11111111";  -- 15E0 = FF
      when "1010111100001" =>  data <= "11111111";  -- 15E1 = FF
      when "1010111100010" =>  data <= "11111111";  -- 15E2 = FF
      when "1010111100011" =>  data <= "11111111";  -- 15E3 = FF
      when "1010111100100" =>  data <= "11111111";  -- 15E4 = FF
      when "1010111100101" =>  data <= "11111111";  -- 15E5 = FF
      when "1010111100110" =>  data <= "11111111";  -- 15E6 = FF
      when "1010111100111" =>  data <= "11111111";  -- 15E7 = FF
      when "1010111101000" =>  data <= "11111111";  -- 15E8 = FF
      when "1010111101001" =>  data <= "11111111";  -- 15E9 = FF
      when "1010111101010" =>  data <= "11111111";  -- 15EA = FF
      when "1010111101011" =>  data <= "11111111";  -- 15EB = FF
      when "1010111101100" =>  data <= "11111111";  -- 15EC = FF
      when "1010111101101" =>  data <= "11111111";  -- 15ED = FF
      when "1010111101110" =>  data <= "11111111";  -- 15EE = FF
      when "1010111101111" =>  data <= "11111111";  -- 15EF = FF
      when "1010111110000" =>  data <= "11111111";  -- 15F0 = FF
      when "1010111110001" =>  data <= "11111111";  -- 15F1 = FF
      when "1010111110010" =>  data <= "11111111";  -- 15F2 = FF
      when "1010111110011" =>  data <= "11111111";  -- 15F3 = FF
      when "1010111110100" =>  data <= "11111111";  -- 15F4 = FF
      when "1010111110101" =>  data <= "11111111";  -- 15F5 = FF
      when "1010111110110" =>  data <= "11111111";  -- 15F6 = FF
      when "1010111110111" =>  data <= "11111111";  -- 15F7 = FF
      when "1010111111000" =>  data <= "11111111";  -- 15F8 = FF
      when "1010111111001" =>  data <= "11111111";  -- 15F9 = FF
      when "1010111111010" =>  data <= "11111111";  -- 15FA = FF
      when "1010111111011" =>  data <= "11111111";  -- 15FB = FF
      when "1010111111100" =>  data <= "11111111";  -- 15FC = FF
      when "1010111111101" =>  data <= "11111111";  -- 15FD = FF
      when "1010111111110" =>  data <= "11111111";  -- 15FE = FF
      when "1010111111111" =>  data <= "11111111";  -- 15FF = FF
      when "1011000000000" =>  data <= "11111111";  -- 1600 = FF
      when "1011000000001" =>  data <= "11111111";  -- 1601 = FF
      when "1011000000010" =>  data <= "11111111";  -- 1602 = FF
      when "1011000000011" =>  data <= "11111111";  -- 1603 = FF
      when "1011000000100" =>  data <= "11111111";  -- 1604 = FF
      when "1011000000101" =>  data <= "11111111";  -- 1605 = FF
      when "1011000000110" =>  data <= "11111111";  -- 1606 = FF
      when "1011000000111" =>  data <= "11111111";  -- 1607 = FF
      when "1011000001000" =>  data <= "11111111";  -- 1608 = FF
      when "1011000001001" =>  data <= "11111111";  -- 1609 = FF
      when "1011000001010" =>  data <= "11111111";  -- 160A = FF
      when "1011000001011" =>  data <= "11111111";  -- 160B = FF
      when "1011000001100" =>  data <= "11111111";  -- 160C = FF
      when "1011000001101" =>  data <= "11111111";  -- 160D = FF
      when "1011000001110" =>  data <= "11111111";  -- 160E = FF
      when "1011000001111" =>  data <= "11111111";  -- 160F = FF
      when "1011000010000" =>  data <= "11111111";  -- 1610 = FF
      when "1011000010001" =>  data <= "11111111";  -- 1611 = FF
      when "1011000010010" =>  data <= "11111111";  -- 1612 = FF
      when "1011000010011" =>  data <= "11111111";  -- 1613 = FF
      when "1011000010100" =>  data <= "11111111";  -- 1614 = FF
      when "1011000010101" =>  data <= "11111111";  -- 1615 = FF
      when "1011000010110" =>  data <= "11111111";  -- 1616 = FF
      when "1011000010111" =>  data <= "11111111";  -- 1617 = FF
      when "1011000011000" =>  data <= "11111111";  -- 1618 = FF
      when "1011000011001" =>  data <= "11111111";  -- 1619 = FF
      when "1011000011010" =>  data <= "11111111";  -- 161A = FF
      when "1011000011011" =>  data <= "11111111";  -- 161B = FF
      when "1011000011100" =>  data <= "11111111";  -- 161C = FF
      when "1011000011101" =>  data <= "11111111";  -- 161D = FF
      when "1011000011110" =>  data <= "11111111";  -- 161E = FF
      when "1011000011111" =>  data <= "11111111";  -- 161F = FF
      when "1011000100000" =>  data <= "11111111";  -- 1620 = FF
      when "1011000100001" =>  data <= "11111111";  -- 1621 = FF
      when "1011000100010" =>  data <= "11111111";  -- 1622 = FF
      when "1011000100011" =>  data <= "11111111";  -- 1623 = FF
      when "1011000100100" =>  data <= "11111111";  -- 1624 = FF
      when "1011000100101" =>  data <= "11111111";  -- 1625 = FF
      when "1011000100110" =>  data <= "11111111";  -- 1626 = FF
      when "1011000100111" =>  data <= "11111111";  -- 1627 = FF
      when "1011000101000" =>  data <= "11111111";  -- 1628 = FF
      when "1011000101001" =>  data <= "11111111";  -- 1629 = FF
      when "1011000101010" =>  data <= "11111111";  -- 162A = FF
      when "1011000101011" =>  data <= "11111111";  -- 162B = FF
      when "1011000101100" =>  data <= "11111111";  -- 162C = FF
      when "1011000101101" =>  data <= "11111111";  -- 162D = FF
      when "1011000101110" =>  data <= "11111111";  -- 162E = FF
      when "1011000101111" =>  data <= "11111111";  -- 162F = FF
      when "1011000110000" =>  data <= "11111111";  -- 1630 = FF
      when "1011000110001" =>  data <= "11111111";  -- 1631 = FF
      when "1011000110010" =>  data <= "11111111";  -- 1632 = FF
      when "1011000110011" =>  data <= "11111111";  -- 1633 = FF
      when "1011000110100" =>  data <= "11111111";  -- 1634 = FF
      when "1011000110101" =>  data <= "11111111";  -- 1635 = FF
      when "1011000110110" =>  data <= "11111111";  -- 1636 = FF
      when "1011000110111" =>  data <= "11111111";  -- 1637 = FF
      when "1011000111000" =>  data <= "11111111";  -- 1638 = FF
      when "1011000111001" =>  data <= "11111111";  -- 1639 = FF
      when "1011000111010" =>  data <= "11111111";  -- 163A = FF
      when "1011000111011" =>  data <= "11111111";  -- 163B = FF
      when "1011000111100" =>  data <= "11111111";  -- 163C = FF
      when "1011000111101" =>  data <= "11111111";  -- 163D = FF
      when "1011000111110" =>  data <= "11111111";  -- 163E = FF
      when "1011000111111" =>  data <= "11111111";  -- 163F = FF
      when "1011001000000" =>  data <= "11111111";  -- 1640 = FF
      when "1011001000001" =>  data <= "11111111";  -- 1641 = FF
      when "1011001000010" =>  data <= "11111111";  -- 1642 = FF
      when "1011001000011" =>  data <= "11111111";  -- 1643 = FF
      when "1011001000100" =>  data <= "11111111";  -- 1644 = FF
      when "1011001000101" =>  data <= "11111111";  -- 1645 = FF
      when "1011001000110" =>  data <= "11111111";  -- 1646 = FF
      when "1011001000111" =>  data <= "11111111";  -- 1647 = FF
      when "1011001001000" =>  data <= "11111111";  -- 1648 = FF
      when "1011001001001" =>  data <= "11111111";  -- 1649 = FF
      when "1011001001010" =>  data <= "11111111";  -- 164A = FF
      when "1011001001011" =>  data <= "11111111";  -- 164B = FF
      when "1011001001100" =>  data <= "11111111";  -- 164C = FF
      when "1011001001101" =>  data <= "11111111";  -- 164D = FF
      when "1011001001110" =>  data <= "11111111";  -- 164E = FF
      when "1011001001111" =>  data <= "11111111";  -- 164F = FF
      when "1011001010000" =>  data <= "11111111";  -- 1650 = FF
      when "1011001010001" =>  data <= "11111111";  -- 1651 = FF
      when "1011001010010" =>  data <= "11111111";  -- 1652 = FF
      when "1011001010011" =>  data <= "11111111";  -- 1653 = FF
      when "1011001010100" =>  data <= "11111111";  -- 1654 = FF
      when "1011001010101" =>  data <= "11111111";  -- 1655 = FF
      when "1011001010110" =>  data <= "11111111";  -- 1656 = FF
      when "1011001010111" =>  data <= "11111111";  -- 1657 = FF
      when "1011001011000" =>  data <= "11111111";  -- 1658 = FF
      when "1011001011001" =>  data <= "11111111";  -- 1659 = FF
      when "1011001011010" =>  data <= "11111111";  -- 165A = FF
      when "1011001011011" =>  data <= "11111111";  -- 165B = FF
      when "1011001011100" =>  data <= "11111111";  -- 165C = FF
      when "1011001011101" =>  data <= "11111111";  -- 165D = FF
      when "1011001011110" =>  data <= "11111111";  -- 165E = FF
      when "1011001011111" =>  data <= "11111111";  -- 165F = FF
      when "1011001100000" =>  data <= "11111111";  -- 1660 = FF
      when "1011001100001" =>  data <= "11111111";  -- 1661 = FF
      when "1011001100010" =>  data <= "11111111";  -- 1662 = FF
      when "1011001100011" =>  data <= "11111111";  -- 1663 = FF
      when "1011001100100" =>  data <= "11111111";  -- 1664 = FF
      when "1011001100101" =>  data <= "11111111";  -- 1665 = FF
      when "1011001100110" =>  data <= "11111111";  -- 1666 = FF
      when "1011001100111" =>  data <= "11111111";  -- 1667 = FF
      when "1011001101000" =>  data <= "11111111";  -- 1668 = FF
      when "1011001101001" =>  data <= "11111111";  -- 1669 = FF
      when "1011001101010" =>  data <= "11111111";  -- 166A = FF
      when "1011001101011" =>  data <= "11111111";  -- 166B = FF
      when "1011001101100" =>  data <= "11111111";  -- 166C = FF
      when "1011001101101" =>  data <= "11111111";  -- 166D = FF
      when "1011001101110" =>  data <= "11111111";  -- 166E = FF
      when "1011001101111" =>  data <= "11111111";  -- 166F = FF
      when "1011001110000" =>  data <= "11111111";  -- 1670 = FF
      when "1011001110001" =>  data <= "11111111";  -- 1671 = FF
      when "1011001110010" =>  data <= "11111111";  -- 1672 = FF
      when "1011001110011" =>  data <= "11111111";  -- 1673 = FF
      when "1011001110100" =>  data <= "11111111";  -- 1674 = FF
      when "1011001110101" =>  data <= "11111111";  -- 1675 = FF
      when "1011001110110" =>  data <= "11111111";  -- 1676 = FF
      when "1011001110111" =>  data <= "11111111";  -- 1677 = FF
      when "1011001111000" =>  data <= "11111111";  -- 1678 = FF
      when "1011001111001" =>  data <= "11111111";  -- 1679 = FF
      when "1011001111010" =>  data <= "11111111";  -- 167A = FF
      when "1011001111011" =>  data <= "11111111";  -- 167B = FF
      when "1011001111100" =>  data <= "11111111";  -- 167C = FF
      when "1011001111101" =>  data <= "11111111";  -- 167D = FF
      when "1011001111110" =>  data <= "11111111";  -- 167E = FF
      when "1011001111111" =>  data <= "11111111";  -- 167F = FF
      when "1011010000000" =>  data <= "11111111";  -- 1680 = FF
      when "1011010000001" =>  data <= "11111111";  -- 1681 = FF
      when "1011010000010" =>  data <= "11111111";  -- 1682 = FF
      when "1011010000011" =>  data <= "11111111";  -- 1683 = FF
      when "1011010000100" =>  data <= "11111111";  -- 1684 = FF
      when "1011010000101" =>  data <= "11111111";  -- 1685 = FF
      when "1011010000110" =>  data <= "11111111";  -- 1686 = FF
      when "1011010000111" =>  data <= "11111111";  -- 1687 = FF
      when "1011010001000" =>  data <= "11111111";  -- 1688 = FF
      when "1011010001001" =>  data <= "11111111";  -- 1689 = FF
      when "1011010001010" =>  data <= "11111111";  -- 168A = FF
      when "1011010001011" =>  data <= "11111111";  -- 168B = FF
      when "1011010001100" =>  data <= "11111111";  -- 168C = FF
      when "1011010001101" =>  data <= "11111111";  -- 168D = FF
      when "1011010001110" =>  data <= "11111111";  -- 168E = FF
      when "1011010001111" =>  data <= "11111111";  -- 168F = FF
      when "1011010010000" =>  data <= "11111111";  -- 1690 = FF
      when "1011010010001" =>  data <= "11111111";  -- 1691 = FF
      when "1011010010010" =>  data <= "11111111";  -- 1692 = FF
      when "1011010010011" =>  data <= "11111111";  -- 1693 = FF
      when "1011010010100" =>  data <= "11111111";  -- 1694 = FF
      when "1011010010101" =>  data <= "11111111";  -- 1695 = FF
      when "1011010010110" =>  data <= "11111111";  -- 1696 = FF
      when "1011010010111" =>  data <= "11111111";  -- 1697 = FF
      when "1011010011000" =>  data <= "11111111";  -- 1698 = FF
      when "1011010011001" =>  data <= "11111111";  -- 1699 = FF
      when "1011010011010" =>  data <= "11111111";  -- 169A = FF
      when "1011010011011" =>  data <= "11111111";  -- 169B = FF
      when "1011010011100" =>  data <= "11111111";  -- 169C = FF
      when "1011010011101" =>  data <= "11111111";  -- 169D = FF
      when "1011010011110" =>  data <= "11111111";  -- 169E = FF
      when "1011010011111" =>  data <= "11111111";  -- 169F = FF
      when "1011010100000" =>  data <= "11111111";  -- 16A0 = FF
      when "1011010100001" =>  data <= "11111111";  -- 16A1 = FF
      when "1011010100010" =>  data <= "11111111";  -- 16A2 = FF
      when "1011010100011" =>  data <= "11111111";  -- 16A3 = FF
      when "1011010100100" =>  data <= "11111111";  -- 16A4 = FF
      when "1011010100101" =>  data <= "11111111";  -- 16A5 = FF
      when "1011010100110" =>  data <= "11111111";  -- 16A6 = FF
      when "1011010100111" =>  data <= "11111111";  -- 16A7 = FF
      when "1011010101000" =>  data <= "11111111";  -- 16A8 = FF
      when "1011010101001" =>  data <= "11111111";  -- 16A9 = FF
      when "1011010101010" =>  data <= "11111111";  -- 16AA = FF
      when "1011010101011" =>  data <= "11111111";  -- 16AB = FF
      when "1011010101100" =>  data <= "11111111";  -- 16AC = FF
      when "1011010101101" =>  data <= "11111111";  -- 16AD = FF
      when "1011010101110" =>  data <= "11111111";  -- 16AE = FF
      when "1011010101111" =>  data <= "11111111";  -- 16AF = FF
      when "1011010110000" =>  data <= "11111111";  -- 16B0 = FF
      when "1011010110001" =>  data <= "11111111";  -- 16B1 = FF
      when "1011010110010" =>  data <= "11111111";  -- 16B2 = FF
      when "1011010110011" =>  data <= "11111111";  -- 16B3 = FF
      when "1011010110100" =>  data <= "11111111";  -- 16B4 = FF
      when "1011010110101" =>  data <= "11111111";  -- 16B5 = FF
      when "1011010110110" =>  data <= "11111111";  -- 16B6 = FF
      when "1011010110111" =>  data <= "11111111";  -- 16B7 = FF
      when "1011010111000" =>  data <= "11111111";  -- 16B8 = FF
      when "1011010111001" =>  data <= "11111111";  -- 16B9 = FF
      when "1011010111010" =>  data <= "11111111";  -- 16BA = FF
      when "1011010111011" =>  data <= "11111111";  -- 16BB = FF
      when "1011010111100" =>  data <= "11111111";  -- 16BC = FF
      when "1011010111101" =>  data <= "11111111";  -- 16BD = FF
      when "1011010111110" =>  data <= "11111111";  -- 16BE = FF
      when "1011010111111" =>  data <= "11111111";  -- 16BF = FF
      when "1011011000000" =>  data <= "11111111";  -- 16C0 = FF
      when "1011011000001" =>  data <= "11111111";  -- 16C1 = FF
      when "1011011000010" =>  data <= "11111111";  -- 16C2 = FF
      when "1011011000011" =>  data <= "11111111";  -- 16C3 = FF
      when "1011011000100" =>  data <= "11111111";  -- 16C4 = FF
      when "1011011000101" =>  data <= "11111111";  -- 16C5 = FF
      when "1011011000110" =>  data <= "11111111";  -- 16C6 = FF
      when "1011011000111" =>  data <= "11111111";  -- 16C7 = FF
      when "1011011001000" =>  data <= "11111111";  -- 16C8 = FF
      when "1011011001001" =>  data <= "11111111";  -- 16C9 = FF
      when "1011011001010" =>  data <= "11111111";  -- 16CA = FF
      when "1011011001011" =>  data <= "11111111";  -- 16CB = FF
      when "1011011001100" =>  data <= "11111111";  -- 16CC = FF
      when "1011011001101" =>  data <= "11111111";  -- 16CD = FF
      when "1011011001110" =>  data <= "11111111";  -- 16CE = FF
      when "1011011001111" =>  data <= "11111111";  -- 16CF = FF
      when "1011011010000" =>  data <= "11111111";  -- 16D0 = FF
      when "1011011010001" =>  data <= "11111111";  -- 16D1 = FF
      when "1011011010010" =>  data <= "11111111";  -- 16D2 = FF
      when "1011011010011" =>  data <= "11111111";  -- 16D3 = FF
      when "1011011010100" =>  data <= "11111111";  -- 16D4 = FF
      when "1011011010101" =>  data <= "11111111";  -- 16D5 = FF
      when "1011011010110" =>  data <= "11111111";  -- 16D6 = FF
      when "1011011010111" =>  data <= "11111111";  -- 16D7 = FF
      when "1011011011000" =>  data <= "11111111";  -- 16D8 = FF
      when "1011011011001" =>  data <= "11111111";  -- 16D9 = FF
      when "1011011011010" =>  data <= "11111111";  -- 16DA = FF
      when "1011011011011" =>  data <= "11111111";  -- 16DB = FF
      when "1011011011100" =>  data <= "11111111";  -- 16DC = FF
      when "1011011011101" =>  data <= "11111111";  -- 16DD = FF
      when "1011011011110" =>  data <= "11111111";  -- 16DE = FF
      when "1011011011111" =>  data <= "11111111";  -- 16DF = FF
      when "1011011100000" =>  data <= "11111111";  -- 16E0 = FF
      when "1011011100001" =>  data <= "11111111";  -- 16E1 = FF
      when "1011011100010" =>  data <= "11111111";  -- 16E2 = FF
      when "1011011100011" =>  data <= "11111111";  -- 16E3 = FF
      when "1011011100100" =>  data <= "11111111";  -- 16E4 = FF
      when "1011011100101" =>  data <= "11111111";  -- 16E5 = FF
      when "1011011100110" =>  data <= "11111111";  -- 16E6 = FF
      when "1011011100111" =>  data <= "11111111";  -- 16E7 = FF
      when "1011011101000" =>  data <= "11111111";  -- 16E8 = FF
      when "1011011101001" =>  data <= "11111111";  -- 16E9 = FF
      when "1011011101010" =>  data <= "11111111";  -- 16EA = FF
      when "1011011101011" =>  data <= "11111111";  -- 16EB = FF
      when "1011011101100" =>  data <= "11111111";  -- 16EC = FF
      when "1011011101101" =>  data <= "11111111";  -- 16ED = FF
      when "1011011101110" =>  data <= "11111111";  -- 16EE = FF
      when "1011011101111" =>  data <= "11111111";  -- 16EF = FF
      when "1011011110000" =>  data <= "11111111";  -- 16F0 = FF
      when "1011011110001" =>  data <= "11111111";  -- 16F1 = FF
      when "1011011110010" =>  data <= "11111111";  -- 16F2 = FF
      when "1011011110011" =>  data <= "11111111";  -- 16F3 = FF
      when "1011011110100" =>  data <= "11111111";  -- 16F4 = FF
      when "1011011110101" =>  data <= "11111111";  -- 16F5 = FF
      when "1011011110110" =>  data <= "11111111";  -- 16F6 = FF
      when "1011011110111" =>  data <= "11111111";  -- 16F7 = FF
      when "1011011111000" =>  data <= "11111111";  -- 16F8 = FF
      when "1011011111001" =>  data <= "11111111";  -- 16F9 = FF
      when "1011011111010" =>  data <= "11111111";  -- 16FA = FF
      when "1011011111011" =>  data <= "11111111";  -- 16FB = FF
      when "1011011111100" =>  data <= "11111111";  -- 16FC = FF
      when "1011011111101" =>  data <= "11111111";  -- 16FD = FF
      when "1011011111110" =>  data <= "11111111";  -- 16FE = FF
      when "1011011111111" =>  data <= "11111111";  -- 16FF = FF
      when "1011100000000" =>  data <= "11111111";  -- 1700 = FF
      when "1011100000001" =>  data <= "11111111";  -- 1701 = FF
      when "1011100000010" =>  data <= "11111111";  -- 1702 = FF
      when "1011100000011" =>  data <= "11111111";  -- 1703 = FF
      when "1011100000100" =>  data <= "11111111";  -- 1704 = FF
      when "1011100000101" =>  data <= "11111111";  -- 1705 = FF
      when "1011100000110" =>  data <= "11111111";  -- 1706 = FF
      when "1011100000111" =>  data <= "11111111";  -- 1707 = FF
      when "1011100001000" =>  data <= "11111111";  -- 1708 = FF
      when "1011100001001" =>  data <= "11111111";  -- 1709 = FF
      when "1011100001010" =>  data <= "11111111";  -- 170A = FF
      when "1011100001011" =>  data <= "11111111";  -- 170B = FF
      when "1011100001100" =>  data <= "11111111";  -- 170C = FF
      when "1011100001101" =>  data <= "11111111";  -- 170D = FF
      when "1011100001110" =>  data <= "11111111";  -- 170E = FF
      when "1011100001111" =>  data <= "11111111";  -- 170F = FF
      when "1011100010000" =>  data <= "11111111";  -- 1710 = FF
      when "1011100010001" =>  data <= "11111111";  -- 1711 = FF
      when "1011100010010" =>  data <= "11111111";  -- 1712 = FF
      when "1011100010011" =>  data <= "11111111";  -- 1713 = FF
      when "1011100010100" =>  data <= "11111111";  -- 1714 = FF
      when "1011100010101" =>  data <= "11111111";  -- 1715 = FF
      when "1011100010110" =>  data <= "11111111";  -- 1716 = FF
      when "1011100010111" =>  data <= "11111111";  -- 1717 = FF
      when "1011100011000" =>  data <= "11111111";  -- 1718 = FF
      when "1011100011001" =>  data <= "11111111";  -- 1719 = FF
      when "1011100011010" =>  data <= "11111111";  -- 171A = FF
      when "1011100011011" =>  data <= "11111111";  -- 171B = FF
      when "1011100011100" =>  data <= "11111111";  -- 171C = FF
      when "1011100011101" =>  data <= "11111111";  -- 171D = FF
      when "1011100011110" =>  data <= "11111111";  -- 171E = FF
      when "1011100011111" =>  data <= "11111111";  -- 171F = FF
      when "1011100100000" =>  data <= "11111111";  -- 1720 = FF
      when "1011100100001" =>  data <= "11111111";  -- 1721 = FF
      when "1011100100010" =>  data <= "11111111";  -- 1722 = FF
      when "1011100100011" =>  data <= "11111111";  -- 1723 = FF
      when "1011100100100" =>  data <= "11111111";  -- 1724 = FF
      when "1011100100101" =>  data <= "11111111";  -- 1725 = FF
      when "1011100100110" =>  data <= "11111111";  -- 1726 = FF
      when "1011100100111" =>  data <= "11111111";  -- 1727 = FF
      when "1011100101000" =>  data <= "11111111";  -- 1728 = FF
      when "1011100101001" =>  data <= "11111111";  -- 1729 = FF
      when "1011100101010" =>  data <= "11111111";  -- 172A = FF
      when "1011100101011" =>  data <= "11111111";  -- 172B = FF
      when "1011100101100" =>  data <= "11111111";  -- 172C = FF
      when "1011100101101" =>  data <= "11111111";  -- 172D = FF
      when "1011100101110" =>  data <= "11111111";  -- 172E = FF
      when "1011100101111" =>  data <= "11111111";  -- 172F = FF
      when "1011100110000" =>  data <= "11111111";  -- 1730 = FF
      when "1011100110001" =>  data <= "11111111";  -- 1731 = FF
      when "1011100110010" =>  data <= "11111111";  -- 1732 = FF
      when "1011100110011" =>  data <= "11111111";  -- 1733 = FF
      when "1011100110100" =>  data <= "11111111";  -- 1734 = FF
      when "1011100110101" =>  data <= "11111111";  -- 1735 = FF
      when "1011100110110" =>  data <= "11111111";  -- 1736 = FF
      when "1011100110111" =>  data <= "11111111";  -- 1737 = FF
      when "1011100111000" =>  data <= "11111111";  -- 1738 = FF
      when "1011100111001" =>  data <= "11111111";  -- 1739 = FF
      when "1011100111010" =>  data <= "11111111";  -- 173A = FF
      when "1011100111011" =>  data <= "11111111";  -- 173B = FF
      when "1011100111100" =>  data <= "11111111";  -- 173C = FF
      when "1011100111101" =>  data <= "11111111";  -- 173D = FF
      when "1011100111110" =>  data <= "11111111";  -- 173E = FF
      when "1011100111111" =>  data <= "11111111";  -- 173F = FF
      when "1011101000000" =>  data <= "11111111";  -- 1740 = FF
      when "1011101000001" =>  data <= "11111111";  -- 1741 = FF
      when "1011101000010" =>  data <= "11111111";  -- 1742 = FF
      when "1011101000011" =>  data <= "11111111";  -- 1743 = FF
      when "1011101000100" =>  data <= "11111111";  -- 1744 = FF
      when "1011101000101" =>  data <= "11111111";  -- 1745 = FF
      when "1011101000110" =>  data <= "11111111";  -- 1746 = FF
      when "1011101000111" =>  data <= "11111111";  -- 1747 = FF
      when "1011101001000" =>  data <= "11111111";  -- 1748 = FF
      when "1011101001001" =>  data <= "11111111";  -- 1749 = FF
      when "1011101001010" =>  data <= "11111111";  -- 174A = FF
      when "1011101001011" =>  data <= "11111111";  -- 174B = FF
      when "1011101001100" =>  data <= "11111111";  -- 174C = FF
      when "1011101001101" =>  data <= "11111111";  -- 174D = FF
      when "1011101001110" =>  data <= "11111111";  -- 174E = FF
      when "1011101001111" =>  data <= "11111111";  -- 174F = FF
      when "1011101010000" =>  data <= "11111111";  -- 1750 = FF
      when "1011101010001" =>  data <= "11111111";  -- 1751 = FF
      when "1011101010010" =>  data <= "11111111";  -- 1752 = FF
      when "1011101010011" =>  data <= "11111111";  -- 1753 = FF
      when "1011101010100" =>  data <= "11111111";  -- 1754 = FF
      when "1011101010101" =>  data <= "11111111";  -- 1755 = FF
      when "1011101010110" =>  data <= "11111111";  -- 1756 = FF
      when "1011101010111" =>  data <= "11111111";  -- 1757 = FF
      when "1011101011000" =>  data <= "11111111";  -- 1758 = FF
      when "1011101011001" =>  data <= "11111111";  -- 1759 = FF
      when "1011101011010" =>  data <= "11111111";  -- 175A = FF
      when "1011101011011" =>  data <= "11111111";  -- 175B = FF
      when "1011101011100" =>  data <= "11111111";  -- 175C = FF
      when "1011101011101" =>  data <= "11111111";  -- 175D = FF
      when "1011101011110" =>  data <= "11111111";  -- 175E = FF
      when "1011101011111" =>  data <= "11111111";  -- 175F = FF
      when "1011101100000" =>  data <= "11111111";  -- 1760 = FF
      when "1011101100001" =>  data <= "11111111";  -- 1761 = FF
      when "1011101100010" =>  data <= "11111111";  -- 1762 = FF
      when "1011101100011" =>  data <= "11111111";  -- 1763 = FF
      when "1011101100100" =>  data <= "11111111";  -- 1764 = FF
      when "1011101100101" =>  data <= "11111111";  -- 1765 = FF
      when "1011101100110" =>  data <= "11111111";  -- 1766 = FF
      when "1011101100111" =>  data <= "11111111";  -- 1767 = FF
      when "1011101101000" =>  data <= "11111111";  -- 1768 = FF
      when "1011101101001" =>  data <= "11111111";  -- 1769 = FF
      when "1011101101010" =>  data <= "11111111";  -- 176A = FF
      when "1011101101011" =>  data <= "11111111";  -- 176B = FF
      when "1011101101100" =>  data <= "11111111";  -- 176C = FF
      when "1011101101101" =>  data <= "11111111";  -- 176D = FF
      when "1011101101110" =>  data <= "11111111";  -- 176E = FF
      when "1011101101111" =>  data <= "11111111";  -- 176F = FF
      when "1011101110000" =>  data <= "11111111";  -- 1770 = FF
      when "1011101110001" =>  data <= "11111111";  -- 1771 = FF
      when "1011101110010" =>  data <= "11111111";  -- 1772 = FF
      when "1011101110011" =>  data <= "11111111";  -- 1773 = FF
      when "1011101110100" =>  data <= "11111111";  -- 1774 = FF
      when "1011101110101" =>  data <= "11111111";  -- 1775 = FF
      when "1011101110110" =>  data <= "11111111";  -- 1776 = FF
      when "1011101110111" =>  data <= "11111111";  -- 1777 = FF
      when "1011101111000" =>  data <= "11111111";  -- 1778 = FF
      when "1011101111001" =>  data <= "11111111";  -- 1779 = FF
      when "1011101111010" =>  data <= "11111111";  -- 177A = FF
      when "1011101111011" =>  data <= "11111111";  -- 177B = FF
      when "1011101111100" =>  data <= "11111111";  -- 177C = FF
      when "1011101111101" =>  data <= "11111111";  -- 177D = FF
      when "1011101111110" =>  data <= "11111111";  -- 177E = FF
      when "1011101111111" =>  data <= "11111111";  -- 177F = FF
      when "1011110000000" =>  data <= "11111111";  -- 1780 = FF
      when "1011110000001" =>  data <= "11111111";  -- 1781 = FF
      when "1011110000010" =>  data <= "11111111";  -- 1782 = FF
      when "1011110000011" =>  data <= "11111111";  -- 1783 = FF
      when "1011110000100" =>  data <= "11111111";  -- 1784 = FF
      when "1011110000101" =>  data <= "11111111";  -- 1785 = FF
      when "1011110000110" =>  data <= "11111111";  -- 1786 = FF
      when "1011110000111" =>  data <= "11111111";  -- 1787 = FF
      when "1011110001000" =>  data <= "11111111";  -- 1788 = FF
      when "1011110001001" =>  data <= "11111111";  -- 1789 = FF
      when "1011110001010" =>  data <= "11111111";  -- 178A = FF
      when "1011110001011" =>  data <= "11111111";  -- 178B = FF
      when "1011110001100" =>  data <= "11111111";  -- 178C = FF
      when "1011110001101" =>  data <= "11111111";  -- 178D = FF
      when "1011110001110" =>  data <= "11111111";  -- 178E = FF
      when "1011110001111" =>  data <= "11111111";  -- 178F = FF
      when "1011110010000" =>  data <= "11111111";  -- 1790 = FF
      when "1011110010001" =>  data <= "11111111";  -- 1791 = FF
      when "1011110010010" =>  data <= "11111111";  -- 1792 = FF
      when "1011110010011" =>  data <= "11111111";  -- 1793 = FF
      when "1011110010100" =>  data <= "11111111";  -- 1794 = FF
      when "1011110010101" =>  data <= "11111111";  -- 1795 = FF
      when "1011110010110" =>  data <= "11111111";  -- 1796 = FF
      when "1011110010111" =>  data <= "11111111";  -- 1797 = FF
      when "1011110011000" =>  data <= "11111111";  -- 1798 = FF
      when "1011110011001" =>  data <= "11111111";  -- 1799 = FF
      when "1011110011010" =>  data <= "11111111";  -- 179A = FF
      when "1011110011011" =>  data <= "11111111";  -- 179B = FF
      when "1011110011100" =>  data <= "11111111";  -- 179C = FF
      when "1011110011101" =>  data <= "11111111";  -- 179D = FF
      when "1011110011110" =>  data <= "11111111";  -- 179E = FF
      when "1011110011111" =>  data <= "11111111";  -- 179F = FF
      when "1011110100000" =>  data <= "11111111";  -- 17A0 = FF
      when "1011110100001" =>  data <= "11111111";  -- 17A1 = FF
      when "1011110100010" =>  data <= "11111111";  -- 17A2 = FF
      when "1011110100011" =>  data <= "11111111";  -- 17A3 = FF
      when "1011110100100" =>  data <= "11111111";  -- 17A4 = FF
      when "1011110100101" =>  data <= "11111111";  -- 17A5 = FF
      when "1011110100110" =>  data <= "11111111";  -- 17A6 = FF
      when "1011110100111" =>  data <= "11111111";  -- 17A7 = FF
      when "1011110101000" =>  data <= "11111111";  -- 17A8 = FF
      when "1011110101001" =>  data <= "11111111";  -- 17A9 = FF
      when "1011110101010" =>  data <= "11111111";  -- 17AA = FF
      when "1011110101011" =>  data <= "11111111";  -- 17AB = FF
      when "1011110101100" =>  data <= "11111111";  -- 17AC = FF
      when "1011110101101" =>  data <= "11111111";  -- 17AD = FF
      when "1011110101110" =>  data <= "11111111";  -- 17AE = FF
      when "1011110101111" =>  data <= "11111111";  -- 17AF = FF
      when "1011110110000" =>  data <= "11111111";  -- 17B0 = FF
      when "1011110110001" =>  data <= "11111111";  -- 17B1 = FF
      when "1011110110010" =>  data <= "11111111";  -- 17B2 = FF
      when "1011110110011" =>  data <= "11111111";  -- 17B3 = FF
      when "1011110110100" =>  data <= "11111111";  -- 17B4 = FF
      when "1011110110101" =>  data <= "11111111";  -- 17B5 = FF
      when "1011110110110" =>  data <= "11111111";  -- 17B6 = FF
      when "1011110110111" =>  data <= "11111111";  -- 17B7 = FF
      when "1011110111000" =>  data <= "11111111";  -- 17B8 = FF
      when "1011110111001" =>  data <= "11111111";  -- 17B9 = FF
      when "1011110111010" =>  data <= "11111111";  -- 17BA = FF
      when "1011110111011" =>  data <= "11111111";  -- 17BB = FF
      when "1011110111100" =>  data <= "11111111";  -- 17BC = FF
      when "1011110111101" =>  data <= "11111111";  -- 17BD = FF
      when "1011110111110" =>  data <= "11111111";  -- 17BE = FF
      when "1011110111111" =>  data <= "11111111";  -- 17BF = FF
      when "1011111000000" =>  data <= "11111111";  -- 17C0 = FF
      when "1011111000001" =>  data <= "11111111";  -- 17C1 = FF
      when "1011111000010" =>  data <= "11111111";  -- 17C2 = FF
      when "1011111000011" =>  data <= "11111111";  -- 17C3 = FF
      when "1011111000100" =>  data <= "11111111";  -- 17C4 = FF
      when "1011111000101" =>  data <= "11111111";  -- 17C5 = FF
      when "1011111000110" =>  data <= "11111111";  -- 17C6 = FF
      when "1011111000111" =>  data <= "11111111";  -- 17C7 = FF
      when "1011111001000" =>  data <= "11111111";  -- 17C8 = FF
      when "1011111001001" =>  data <= "11111111";  -- 17C9 = FF
      when "1011111001010" =>  data <= "11111111";  -- 17CA = FF
      when "1011111001011" =>  data <= "11111111";  -- 17CB = FF
      when "1011111001100" =>  data <= "11111111";  -- 17CC = FF
      when "1011111001101" =>  data <= "11111111";  -- 17CD = FF
      when "1011111001110" =>  data <= "11111111";  -- 17CE = FF
      when "1011111001111" =>  data <= "11111111";  -- 17CF = FF
      when "1011111010000" =>  data <= "11111111";  -- 17D0 = FF
      when "1011111010001" =>  data <= "11111111";  -- 17D1 = FF
      when "1011111010010" =>  data <= "11111111";  -- 17D2 = FF
      when "1011111010011" =>  data <= "11111111";  -- 17D3 = FF
      when "1011111010100" =>  data <= "11111111";  -- 17D4 = FF
      when "1011111010101" =>  data <= "11111111";  -- 17D5 = FF
      when "1011111010110" =>  data <= "11111111";  -- 17D6 = FF
      when "1011111010111" =>  data <= "11111111";  -- 17D7 = FF
      when "1011111011000" =>  data <= "11111111";  -- 17D8 = FF
      when "1011111011001" =>  data <= "11111111";  -- 17D9 = FF
      when "1011111011010" =>  data <= "11111111";  -- 17DA = FF
      when "1011111011011" =>  data <= "11111111";  -- 17DB = FF
      when "1011111011100" =>  data <= "11111111";  -- 17DC = FF
      when "1011111011101" =>  data <= "11111111";  -- 17DD = FF
      when "1011111011110" =>  data <= "11111111";  -- 17DE = FF
      when "1011111011111" =>  data <= "11111111";  -- 17DF = FF
      when "1011111100000" =>  data <= "11111111";  -- 17E0 = FF
      when "1011111100001" =>  data <= "11111111";  -- 17E1 = FF
      when "1011111100010" =>  data <= "11111111";  -- 17E2 = FF
      when "1011111100011" =>  data <= "11111111";  -- 17E3 = FF
      when "1011111100100" =>  data <= "11111111";  -- 17E4 = FF
      when "1011111100101" =>  data <= "11111111";  -- 17E5 = FF
      when "1011111100110" =>  data <= "11111111";  -- 17E6 = FF
      when "1011111100111" =>  data <= "11111111";  -- 17E7 = FF
      when "1011111101000" =>  data <= "11111111";  -- 17E8 = FF
      when "1011111101001" =>  data <= "11111111";  -- 17E9 = FF
      when "1011111101010" =>  data <= "11111111";  -- 17EA = FF
      when "1011111101011" =>  data <= "11111111";  -- 17EB = FF
      when "1011111101100" =>  data <= "11111111";  -- 17EC = FF
      when "1011111101101" =>  data <= "11111111";  -- 17ED = FF
      when "1011111101110" =>  data <= "11111111";  -- 17EE = FF
      when "1011111101111" =>  data <= "11111111";  -- 17EF = FF
      when "1011111110000" =>  data <= "11111111";  -- 17F0 = FF
      when "1011111110001" =>  data <= "11111111";  -- 17F1 = FF
      when "1011111110010" =>  data <= "11111111";  -- 17F2 = FF
      when "1011111110011" =>  data <= "11111111";  -- 17F3 = FF
      when "1011111110100" =>  data <= "11111111";  -- 17F4 = FF
      when "1011111110101" =>  data <= "11111111";  -- 17F5 = FF
      when "1011111110110" =>  data <= "11111111";  -- 17F6 = FF
      when "1011111110111" =>  data <= "11111111";  -- 17F7 = FF
      when "1011111111000" =>  data <= "11111111";  -- 17F8 = FF
      when "1011111111001" =>  data <= "11111111";  -- 17F9 = FF
      when "1011111111010" =>  data <= "11111111";  -- 17FA = FF
      when "1011111111011" =>  data <= "11111111";  -- 17FB = FF
      when "1011111111100" =>  data <= "11111111";  -- 17FC = FF
      when "1011111111101" =>  data <= "11111111";  -- 17FD = FF
      when "1011111111110" =>  data <= "11111111";  -- 17FE = FF
      when "1011111111111" =>  data <= "11111111";  -- 17FF = FF
      when "1100000000000" =>  data <= "11111111";  -- 1800 = FF
      when "1100000000001" =>  data <= "11111111";  -- 1801 = FF
      when "1100000000010" =>  data <= "11111111";  -- 1802 = FF
      when "1100000000011" =>  data <= "11111111";  -- 1803 = FF
      when "1100000000100" =>  data <= "11111111";  -- 1804 = FF
      when "1100000000101" =>  data <= "11111111";  -- 1805 = FF
      when "1100000000110" =>  data <= "11111111";  -- 1806 = FF
      when "1100000000111" =>  data <= "11111111";  -- 1807 = FF
      when "1100000001000" =>  data <= "11111111";  -- 1808 = FF
      when "1100000001001" =>  data <= "11111111";  -- 1809 = FF
      when "1100000001010" =>  data <= "11111111";  -- 180A = FF
      when "1100000001011" =>  data <= "11111111";  -- 180B = FF
      when "1100000001100" =>  data <= "11111111";  -- 180C = FF
      when "1100000001101" =>  data <= "11111111";  -- 180D = FF
      when "1100000001110" =>  data <= "11111111";  -- 180E = FF
      when "1100000001111" =>  data <= "11111111";  -- 180F = FF
      when "1100000010000" =>  data <= "11111111";  -- 1810 = FF
      when "1100000010001" =>  data <= "11111111";  -- 1811 = FF
      when "1100000010010" =>  data <= "11111111";  -- 1812 = FF
      when "1100000010011" =>  data <= "11111111";  -- 1813 = FF
      when "1100000010100" =>  data <= "11111111";  -- 1814 = FF
      when "1100000010101" =>  data <= "11111111";  -- 1815 = FF
      when "1100000010110" =>  data <= "11111111";  -- 1816 = FF
      when "1100000010111" =>  data <= "11111111";  -- 1817 = FF
      when "1100000011000" =>  data <= "11111111";  -- 1818 = FF
      when "1100000011001" =>  data <= "11111111";  -- 1819 = FF
      when "1100000011010" =>  data <= "11111111";  -- 181A = FF
      when "1100000011011" =>  data <= "11111111";  -- 181B = FF
      when "1100000011100" =>  data <= "11111111";  -- 181C = FF
      when "1100000011101" =>  data <= "11111111";  -- 181D = FF
      when "1100000011110" =>  data <= "11111111";  -- 181E = FF
      when "1100000011111" =>  data <= "11111111";  -- 181F = FF
      when "1100000100000" =>  data <= "11111111";  -- 1820 = FF
      when "1100000100001" =>  data <= "11111111";  -- 1821 = FF
      when "1100000100010" =>  data <= "11111111";  -- 1822 = FF
      when "1100000100011" =>  data <= "11111111";  -- 1823 = FF
      when "1100000100100" =>  data <= "11111111";  -- 1824 = FF
      when "1100000100101" =>  data <= "11111111";  -- 1825 = FF
      when "1100000100110" =>  data <= "11111111";  -- 1826 = FF
      when "1100000100111" =>  data <= "11111111";  -- 1827 = FF
      when "1100000101000" =>  data <= "11111111";  -- 1828 = FF
      when "1100000101001" =>  data <= "11111111";  -- 1829 = FF
      when "1100000101010" =>  data <= "11111111";  -- 182A = FF
      when "1100000101011" =>  data <= "11111111";  -- 182B = FF
      when "1100000101100" =>  data <= "11111111";  -- 182C = FF
      when "1100000101101" =>  data <= "11111111";  -- 182D = FF
      when "1100000101110" =>  data <= "11111111";  -- 182E = FF
      when "1100000101111" =>  data <= "11111111";  -- 182F = FF
      when "1100000110000" =>  data <= "11111111";  -- 1830 = FF
      when "1100000110001" =>  data <= "11111111";  -- 1831 = FF
      when "1100000110010" =>  data <= "11111111";  -- 1832 = FF
      when "1100000110011" =>  data <= "11111111";  -- 1833 = FF
      when "1100000110100" =>  data <= "11111111";  -- 1834 = FF
      when "1100000110101" =>  data <= "11111111";  -- 1835 = FF
      when "1100000110110" =>  data <= "11111111";  -- 1836 = FF
      when "1100000110111" =>  data <= "11111111";  -- 1837 = FF
      when "1100000111000" =>  data <= "11111111";  -- 1838 = FF
      when "1100000111001" =>  data <= "11111111";  -- 1839 = FF
      when "1100000111010" =>  data <= "11111111";  -- 183A = FF
      when "1100000111011" =>  data <= "11111111";  -- 183B = FF
      when "1100000111100" =>  data <= "11111111";  -- 183C = FF
      when "1100000111101" =>  data <= "11111111";  -- 183D = FF
      when "1100000111110" =>  data <= "11111111";  -- 183E = FF
      when "1100000111111" =>  data <= "11111111";  -- 183F = FF
      when "1100001000000" =>  data <= "11111111";  -- 1840 = FF
      when "1100001000001" =>  data <= "11111111";  -- 1841 = FF
      when "1100001000010" =>  data <= "11111111";  -- 1842 = FF
      when "1100001000011" =>  data <= "11111111";  -- 1843 = FF
      when "1100001000100" =>  data <= "11111111";  -- 1844 = FF
      when "1100001000101" =>  data <= "11111111";  -- 1845 = FF
      when "1100001000110" =>  data <= "11111111";  -- 1846 = FF
      when "1100001000111" =>  data <= "11111111";  -- 1847 = FF
      when "1100001001000" =>  data <= "11111111";  -- 1848 = FF
      when "1100001001001" =>  data <= "11111111";  -- 1849 = FF
      when "1100001001010" =>  data <= "11111111";  -- 184A = FF
      when "1100001001011" =>  data <= "11111111";  -- 184B = FF
      when "1100001001100" =>  data <= "11111111";  -- 184C = FF
      when "1100001001101" =>  data <= "11111111";  -- 184D = FF
      when "1100001001110" =>  data <= "11111111";  -- 184E = FF
      when "1100001001111" =>  data <= "11111111";  -- 184F = FF
      when "1100001010000" =>  data <= "11111111";  -- 1850 = FF
      when "1100001010001" =>  data <= "11111111";  -- 1851 = FF
      when "1100001010010" =>  data <= "11111111";  -- 1852 = FF
      when "1100001010011" =>  data <= "11111111";  -- 1853 = FF
      when "1100001010100" =>  data <= "11111111";  -- 1854 = FF
      when "1100001010101" =>  data <= "11111111";  -- 1855 = FF
      when "1100001010110" =>  data <= "11111111";  -- 1856 = FF
      when "1100001010111" =>  data <= "11111111";  -- 1857 = FF
      when "1100001011000" =>  data <= "11111111";  -- 1858 = FF
      when "1100001011001" =>  data <= "11111111";  -- 1859 = FF
      when "1100001011010" =>  data <= "11111111";  -- 185A = FF
      when "1100001011011" =>  data <= "11111111";  -- 185B = FF
      when "1100001011100" =>  data <= "11111111";  -- 185C = FF
      when "1100001011101" =>  data <= "11111111";  -- 185D = FF
      when "1100001011110" =>  data <= "11111111";  -- 185E = FF
      when "1100001011111" =>  data <= "11111111";  -- 185F = FF
      when "1100001100000" =>  data <= "11111111";  -- 1860 = FF
      when "1100001100001" =>  data <= "11111111";  -- 1861 = FF
      when "1100001100010" =>  data <= "11111111";  -- 1862 = FF
      when "1100001100011" =>  data <= "11111111";  -- 1863 = FF
      when "1100001100100" =>  data <= "11111111";  -- 1864 = FF
      when "1100001100101" =>  data <= "11111111";  -- 1865 = FF
      when "1100001100110" =>  data <= "11111111";  -- 1866 = FF
      when "1100001100111" =>  data <= "11111111";  -- 1867 = FF
      when "1100001101000" =>  data <= "11111111";  -- 1868 = FF
      when "1100001101001" =>  data <= "11111111";  -- 1869 = FF
      when "1100001101010" =>  data <= "11111111";  -- 186A = FF
      when "1100001101011" =>  data <= "11111111";  -- 186B = FF
      when "1100001101100" =>  data <= "11111111";  -- 186C = FF
      when "1100001101101" =>  data <= "11111111";  -- 186D = FF
      when "1100001101110" =>  data <= "11111111";  -- 186E = FF
      when "1100001101111" =>  data <= "11111111";  -- 186F = FF
      when "1100001110000" =>  data <= "11111111";  -- 1870 = FF
      when "1100001110001" =>  data <= "11111111";  -- 1871 = FF
      when "1100001110010" =>  data <= "11111111";  -- 1872 = FF
      when "1100001110011" =>  data <= "11111111";  -- 1873 = FF
      when "1100001110100" =>  data <= "11111111";  -- 1874 = FF
      when "1100001110101" =>  data <= "11111111";  -- 1875 = FF
      when "1100001110110" =>  data <= "11111111";  -- 1876 = FF
      when "1100001110111" =>  data <= "11111111";  -- 1877 = FF
      when "1100001111000" =>  data <= "11111111";  -- 1878 = FF
      when "1100001111001" =>  data <= "11111111";  -- 1879 = FF
      when "1100001111010" =>  data <= "11111111";  -- 187A = FF
      when "1100001111011" =>  data <= "11111111";  -- 187B = FF
      when "1100001111100" =>  data <= "11111111";  -- 187C = FF
      when "1100001111101" =>  data <= "11111111";  -- 187D = FF
      when "1100001111110" =>  data <= "11111111";  -- 187E = FF
      when "1100001111111" =>  data <= "11111111";  -- 187F = FF
      when "1100010000000" =>  data <= "11111111";  -- 1880 = FF
      when "1100010000001" =>  data <= "11111111";  -- 1881 = FF
      when "1100010000010" =>  data <= "11111111";  -- 1882 = FF
      when "1100010000011" =>  data <= "11111111";  -- 1883 = FF
      when "1100010000100" =>  data <= "11111111";  -- 1884 = FF
      when "1100010000101" =>  data <= "11111111";  -- 1885 = FF
      when "1100010000110" =>  data <= "11111111";  -- 1886 = FF
      when "1100010000111" =>  data <= "11111111";  -- 1887 = FF
      when "1100010001000" =>  data <= "11111111";  -- 1888 = FF
      when "1100010001001" =>  data <= "11111111";  -- 1889 = FF
      when "1100010001010" =>  data <= "11111111";  -- 188A = FF
      when "1100010001011" =>  data <= "11111111";  -- 188B = FF
      when "1100010001100" =>  data <= "11111111";  -- 188C = FF
      when "1100010001101" =>  data <= "11111111";  -- 188D = FF
      when "1100010001110" =>  data <= "11111111";  -- 188E = FF
      when "1100010001111" =>  data <= "11111111";  -- 188F = FF
      when "1100010010000" =>  data <= "11111111";  -- 1890 = FF
      when "1100010010001" =>  data <= "11111111";  -- 1891 = FF
      when "1100010010010" =>  data <= "11111111";  -- 1892 = FF
      when "1100010010011" =>  data <= "11111111";  -- 1893 = FF
      when "1100010010100" =>  data <= "11111111";  -- 1894 = FF
      when "1100010010101" =>  data <= "11111111";  -- 1895 = FF
      when "1100010010110" =>  data <= "11111111";  -- 1896 = FF
      when "1100010010111" =>  data <= "11111111";  -- 1897 = FF
      when "1100010011000" =>  data <= "11111111";  -- 1898 = FF
      when "1100010011001" =>  data <= "11111111";  -- 1899 = FF
      when "1100010011010" =>  data <= "11111111";  -- 189A = FF
      when "1100010011011" =>  data <= "11111111";  -- 189B = FF
      when "1100010011100" =>  data <= "11111111";  -- 189C = FF
      when "1100010011101" =>  data <= "11111111";  -- 189D = FF
      when "1100010011110" =>  data <= "11111111";  -- 189E = FF
      when "1100010011111" =>  data <= "11111111";  -- 189F = FF
      when "1100010100000" =>  data <= "11111111";  -- 18A0 = FF
      when "1100010100001" =>  data <= "11111111";  -- 18A1 = FF
      when "1100010100010" =>  data <= "11111111";  -- 18A2 = FF
      when "1100010100011" =>  data <= "11111111";  -- 18A3 = FF
      when "1100010100100" =>  data <= "11111111";  -- 18A4 = FF
      when "1100010100101" =>  data <= "11111111";  -- 18A5 = FF
      when "1100010100110" =>  data <= "11111111";  -- 18A6 = FF
      when "1100010100111" =>  data <= "11111111";  -- 18A7 = FF
      when "1100010101000" =>  data <= "11111111";  -- 18A8 = FF
      when "1100010101001" =>  data <= "11111111";  -- 18A9 = FF
      when "1100010101010" =>  data <= "11111111";  -- 18AA = FF
      when "1100010101011" =>  data <= "11111111";  -- 18AB = FF
      when "1100010101100" =>  data <= "11111111";  -- 18AC = FF
      when "1100010101101" =>  data <= "11111111";  -- 18AD = FF
      when "1100010101110" =>  data <= "11111111";  -- 18AE = FF
      when "1100010101111" =>  data <= "11111111";  -- 18AF = FF
      when "1100010110000" =>  data <= "11111111";  -- 18B0 = FF
      when "1100010110001" =>  data <= "11111111";  -- 18B1 = FF
      when "1100010110010" =>  data <= "11111111";  -- 18B2 = FF
      when "1100010110011" =>  data <= "11111111";  -- 18B3 = FF
      when "1100010110100" =>  data <= "11111111";  -- 18B4 = FF
      when "1100010110101" =>  data <= "11111111";  -- 18B5 = FF
      when "1100010110110" =>  data <= "11111111";  -- 18B6 = FF
      when "1100010110111" =>  data <= "11111111";  -- 18B7 = FF
      when "1100010111000" =>  data <= "11111111";  -- 18B8 = FF
      when "1100010111001" =>  data <= "11111111";  -- 18B9 = FF
      when "1100010111010" =>  data <= "11111111";  -- 18BA = FF
      when "1100010111011" =>  data <= "11111111";  -- 18BB = FF
      when "1100010111100" =>  data <= "11111111";  -- 18BC = FF
      when "1100010111101" =>  data <= "11111111";  -- 18BD = FF
      when "1100010111110" =>  data <= "11111111";  -- 18BE = FF
      when "1100010111111" =>  data <= "11111111";  -- 18BF = FF
      when "1100011000000" =>  data <= "11111111";  -- 18C0 = FF
      when "1100011000001" =>  data <= "11111111";  -- 18C1 = FF
      when "1100011000010" =>  data <= "11111111";  -- 18C2 = FF
      when "1100011000011" =>  data <= "11111111";  -- 18C3 = FF
      when "1100011000100" =>  data <= "11111111";  -- 18C4 = FF
      when "1100011000101" =>  data <= "11111111";  -- 18C5 = FF
      when "1100011000110" =>  data <= "11111111";  -- 18C6 = FF
      when "1100011000111" =>  data <= "11111111";  -- 18C7 = FF
      when "1100011001000" =>  data <= "11111111";  -- 18C8 = FF
      when "1100011001001" =>  data <= "11111111";  -- 18C9 = FF
      when "1100011001010" =>  data <= "11111111";  -- 18CA = FF
      when "1100011001011" =>  data <= "11111111";  -- 18CB = FF
      when "1100011001100" =>  data <= "11111111";  -- 18CC = FF
      when "1100011001101" =>  data <= "11111111";  -- 18CD = FF
      when "1100011001110" =>  data <= "11111111";  -- 18CE = FF
      when "1100011001111" =>  data <= "11111111";  -- 18CF = FF
      when "1100011010000" =>  data <= "11111111";  -- 18D0 = FF
      when "1100011010001" =>  data <= "11111111";  -- 18D1 = FF
      when "1100011010010" =>  data <= "11111111";  -- 18D2 = FF
      when "1100011010011" =>  data <= "11111111";  -- 18D3 = FF
      when "1100011010100" =>  data <= "11111111";  -- 18D4 = FF
      when "1100011010101" =>  data <= "11111111";  -- 18D5 = FF
      when "1100011010110" =>  data <= "11111111";  -- 18D6 = FF
      when "1100011010111" =>  data <= "11111111";  -- 18D7 = FF
      when "1100011011000" =>  data <= "11111111";  -- 18D8 = FF
      when "1100011011001" =>  data <= "11111111";  -- 18D9 = FF
      when "1100011011010" =>  data <= "11111111";  -- 18DA = FF
      when "1100011011011" =>  data <= "11111111";  -- 18DB = FF
      when "1100011011100" =>  data <= "11111111";  -- 18DC = FF
      when "1100011011101" =>  data <= "11111111";  -- 18DD = FF
      when "1100011011110" =>  data <= "11111111";  -- 18DE = FF
      when "1100011011111" =>  data <= "11111111";  -- 18DF = FF
      when "1100011100000" =>  data <= "11111111";  -- 18E0 = FF
      when "1100011100001" =>  data <= "11111111";  -- 18E1 = FF
      when "1100011100010" =>  data <= "11111111";  -- 18E2 = FF
      when "1100011100011" =>  data <= "11111111";  -- 18E3 = FF
      when "1100011100100" =>  data <= "11111111";  -- 18E4 = FF
      when "1100011100101" =>  data <= "11111111";  -- 18E5 = FF
      when "1100011100110" =>  data <= "11111111";  -- 18E6 = FF
      when "1100011100111" =>  data <= "11111111";  -- 18E7 = FF
      when "1100011101000" =>  data <= "11111111";  -- 18E8 = FF
      when "1100011101001" =>  data <= "11111111";  -- 18E9 = FF
      when "1100011101010" =>  data <= "11111111";  -- 18EA = FF
      when "1100011101011" =>  data <= "11111111";  -- 18EB = FF
      when "1100011101100" =>  data <= "11111111";  -- 18EC = FF
      when "1100011101101" =>  data <= "11111111";  -- 18ED = FF
      when "1100011101110" =>  data <= "11111111";  -- 18EE = FF
      when "1100011101111" =>  data <= "11111111";  -- 18EF = FF
      when "1100011110000" =>  data <= "11111111";  -- 18F0 = FF
      when "1100011110001" =>  data <= "11111111";  -- 18F1 = FF
      when "1100011110010" =>  data <= "11111111";  -- 18F2 = FF
      when "1100011110011" =>  data <= "11111111";  -- 18F3 = FF
      when "1100011110100" =>  data <= "11111111";  -- 18F4 = FF
      when "1100011110101" =>  data <= "11111111";  -- 18F5 = FF
      when "1100011110110" =>  data <= "11111111";  -- 18F6 = FF
      when "1100011110111" =>  data <= "11111111";  -- 18F7 = FF
      when "1100011111000" =>  data <= "11111111";  -- 18F8 = FF
      when "1100011111001" =>  data <= "11111111";  -- 18F9 = FF
      when "1100011111010" =>  data <= "11111111";  -- 18FA = FF
      when "1100011111011" =>  data <= "11111111";  -- 18FB = FF
      when "1100011111100" =>  data <= "11111111";  -- 18FC = FF
      when "1100011111101" =>  data <= "11111111";  -- 18FD = FF
      when "1100011111110" =>  data <= "11111111";  -- 18FE = FF
      when "1100011111111" =>  data <= "11111111";  -- 18FF = FF
      when "1100100000000" =>  data <= "11111111";  -- 1900 = FF
      when "1100100000001" =>  data <= "11111111";  -- 1901 = FF
      when "1100100000010" =>  data <= "11111111";  -- 1902 = FF
      when "1100100000011" =>  data <= "11111111";  -- 1903 = FF
      when "1100100000100" =>  data <= "11111111";  -- 1904 = FF
      when "1100100000101" =>  data <= "11111111";  -- 1905 = FF
      when "1100100000110" =>  data <= "11111111";  -- 1906 = FF
      when "1100100000111" =>  data <= "11111111";  -- 1907 = FF
      when "1100100001000" =>  data <= "11111111";  -- 1908 = FF
      when "1100100001001" =>  data <= "11111111";  -- 1909 = FF
      when "1100100001010" =>  data <= "11111111";  -- 190A = FF
      when "1100100001011" =>  data <= "11111111";  -- 190B = FF
      when "1100100001100" =>  data <= "11111111";  -- 190C = FF
      when "1100100001101" =>  data <= "11111111";  -- 190D = FF
      when "1100100001110" =>  data <= "11111111";  -- 190E = FF
      when "1100100001111" =>  data <= "11111111";  -- 190F = FF
      when "1100100010000" =>  data <= "11111111";  -- 1910 = FF
      when "1100100010001" =>  data <= "11111111";  -- 1911 = FF
      when "1100100010010" =>  data <= "11111111";  -- 1912 = FF
      when "1100100010011" =>  data <= "11111111";  -- 1913 = FF
      when "1100100010100" =>  data <= "11111111";  -- 1914 = FF
      when "1100100010101" =>  data <= "11111111";  -- 1915 = FF
      when "1100100010110" =>  data <= "11111111";  -- 1916 = FF
      when "1100100010111" =>  data <= "11111111";  -- 1917 = FF
      when "1100100011000" =>  data <= "11111111";  -- 1918 = FF
      when "1100100011001" =>  data <= "11111111";  -- 1919 = FF
      when "1100100011010" =>  data <= "11111111";  -- 191A = FF
      when "1100100011011" =>  data <= "11111111";  -- 191B = FF
      when "1100100011100" =>  data <= "11111111";  -- 191C = FF
      when "1100100011101" =>  data <= "11111111";  -- 191D = FF
      when "1100100011110" =>  data <= "11111111";  -- 191E = FF
      when "1100100011111" =>  data <= "11111111";  -- 191F = FF
      when "1100100100000" =>  data <= "11111111";  -- 1920 = FF
      when "1100100100001" =>  data <= "11111111";  -- 1921 = FF
      when "1100100100010" =>  data <= "11111111";  -- 1922 = FF
      when "1100100100011" =>  data <= "11111111";  -- 1923 = FF
      when "1100100100100" =>  data <= "11111111";  -- 1924 = FF
      when "1100100100101" =>  data <= "11111111";  -- 1925 = FF
      when "1100100100110" =>  data <= "11111111";  -- 1926 = FF
      when "1100100100111" =>  data <= "11111111";  -- 1927 = FF
      when "1100100101000" =>  data <= "11111111";  -- 1928 = FF
      when "1100100101001" =>  data <= "11111111";  -- 1929 = FF
      when "1100100101010" =>  data <= "11111111";  -- 192A = FF
      when "1100100101011" =>  data <= "11111111";  -- 192B = FF
      when "1100100101100" =>  data <= "11111111";  -- 192C = FF
      when "1100100101101" =>  data <= "11111111";  -- 192D = FF
      when "1100100101110" =>  data <= "11111111";  -- 192E = FF
      when "1100100101111" =>  data <= "11111111";  -- 192F = FF
      when "1100100110000" =>  data <= "11111111";  -- 1930 = FF
      when "1100100110001" =>  data <= "11111111";  -- 1931 = FF
      when "1100100110010" =>  data <= "11111111";  -- 1932 = FF
      when "1100100110011" =>  data <= "11111111";  -- 1933 = FF
      when "1100100110100" =>  data <= "11111111";  -- 1934 = FF
      when "1100100110101" =>  data <= "11111111";  -- 1935 = FF
      when "1100100110110" =>  data <= "11111111";  -- 1936 = FF
      when "1100100110111" =>  data <= "11111111";  -- 1937 = FF
      when "1100100111000" =>  data <= "11111111";  -- 1938 = FF
      when "1100100111001" =>  data <= "11111111";  -- 1939 = FF
      when "1100100111010" =>  data <= "11111111";  -- 193A = FF
      when "1100100111011" =>  data <= "11111111";  -- 193B = FF
      when "1100100111100" =>  data <= "11111111";  -- 193C = FF
      when "1100100111101" =>  data <= "11111111";  -- 193D = FF
      when "1100100111110" =>  data <= "11111111";  -- 193E = FF
      when "1100100111111" =>  data <= "11111111";  -- 193F = FF
      when "1100101000000" =>  data <= "11111111";  -- 1940 = FF
      when "1100101000001" =>  data <= "11111111";  -- 1941 = FF
      when "1100101000010" =>  data <= "11111111";  -- 1942 = FF
      when "1100101000011" =>  data <= "11111111";  -- 1943 = FF
      when "1100101000100" =>  data <= "11111111";  -- 1944 = FF
      when "1100101000101" =>  data <= "11111111";  -- 1945 = FF
      when "1100101000110" =>  data <= "11111111";  -- 1946 = FF
      when "1100101000111" =>  data <= "11111111";  -- 1947 = FF
      when "1100101001000" =>  data <= "11111111";  -- 1948 = FF
      when "1100101001001" =>  data <= "11111111";  -- 1949 = FF
      when "1100101001010" =>  data <= "11111111";  -- 194A = FF
      when "1100101001011" =>  data <= "11111111";  -- 194B = FF
      when "1100101001100" =>  data <= "11111111";  -- 194C = FF
      when "1100101001101" =>  data <= "11111111";  -- 194D = FF
      when "1100101001110" =>  data <= "11111111";  -- 194E = FF
      when "1100101001111" =>  data <= "11111111";  -- 194F = FF
      when "1100101010000" =>  data <= "11111111";  -- 1950 = FF
      when "1100101010001" =>  data <= "11111111";  -- 1951 = FF
      when "1100101010010" =>  data <= "11111111";  -- 1952 = FF
      when "1100101010011" =>  data <= "11111111";  -- 1953 = FF
      when "1100101010100" =>  data <= "11111111";  -- 1954 = FF
      when "1100101010101" =>  data <= "11111111";  -- 1955 = FF
      when "1100101010110" =>  data <= "11111111";  -- 1956 = FF
      when "1100101010111" =>  data <= "11111111";  -- 1957 = FF
      when "1100101011000" =>  data <= "11111111";  -- 1958 = FF
      when "1100101011001" =>  data <= "11111111";  -- 1959 = FF
      when "1100101011010" =>  data <= "11111111";  -- 195A = FF
      when "1100101011011" =>  data <= "11111111";  -- 195B = FF
      when "1100101011100" =>  data <= "11111111";  -- 195C = FF
      when "1100101011101" =>  data <= "11111111";  -- 195D = FF
      when "1100101011110" =>  data <= "11111111";  -- 195E = FF
      when "1100101011111" =>  data <= "11111111";  -- 195F = FF
      when "1100101100000" =>  data <= "11111111";  -- 1960 = FF
      when "1100101100001" =>  data <= "11111111";  -- 1961 = FF
      when "1100101100010" =>  data <= "11111111";  -- 1962 = FF
      when "1100101100011" =>  data <= "11111111";  -- 1963 = FF
      when "1100101100100" =>  data <= "11111111";  -- 1964 = FF
      when "1100101100101" =>  data <= "11111111";  -- 1965 = FF
      when "1100101100110" =>  data <= "11111111";  -- 1966 = FF
      when "1100101100111" =>  data <= "11111111";  -- 1967 = FF
      when "1100101101000" =>  data <= "11111111";  -- 1968 = FF
      when "1100101101001" =>  data <= "11111111";  -- 1969 = FF
      when "1100101101010" =>  data <= "11111111";  -- 196A = FF
      when "1100101101011" =>  data <= "11111111";  -- 196B = FF
      when "1100101101100" =>  data <= "11111111";  -- 196C = FF
      when "1100101101101" =>  data <= "11111111";  -- 196D = FF
      when "1100101101110" =>  data <= "11111111";  -- 196E = FF
      when "1100101101111" =>  data <= "11111111";  -- 196F = FF
      when "1100101110000" =>  data <= "11111111";  -- 1970 = FF
      when "1100101110001" =>  data <= "11111111";  -- 1971 = FF
      when "1100101110010" =>  data <= "11111111";  -- 1972 = FF
      when "1100101110011" =>  data <= "11111111";  -- 1973 = FF
      when "1100101110100" =>  data <= "11111111";  -- 1974 = FF
      when "1100101110101" =>  data <= "11111111";  -- 1975 = FF
      when "1100101110110" =>  data <= "11111111";  -- 1976 = FF
      when "1100101110111" =>  data <= "11111111";  -- 1977 = FF
      when "1100101111000" =>  data <= "11111111";  -- 1978 = FF
      when "1100101111001" =>  data <= "11111111";  -- 1979 = FF
      when "1100101111010" =>  data <= "11111111";  -- 197A = FF
      when "1100101111011" =>  data <= "11111111";  -- 197B = FF
      when "1100101111100" =>  data <= "11111111";  -- 197C = FF
      when "1100101111101" =>  data <= "11111111";  -- 197D = FF
      when "1100101111110" =>  data <= "11111111";  -- 197E = FF
      when "1100101111111" =>  data <= "11111111";  -- 197F = FF
      when "1100110000000" =>  data <= "11111111";  -- 1980 = FF
      when "1100110000001" =>  data <= "11111111";  -- 1981 = FF
      when "1100110000010" =>  data <= "11111111";  -- 1982 = FF
      when "1100110000011" =>  data <= "11111111";  -- 1983 = FF
      when "1100110000100" =>  data <= "11111111";  -- 1984 = FF
      when "1100110000101" =>  data <= "11111111";  -- 1985 = FF
      when "1100110000110" =>  data <= "11111111";  -- 1986 = FF
      when "1100110000111" =>  data <= "11111111";  -- 1987 = FF
      when "1100110001000" =>  data <= "11111111";  -- 1988 = FF
      when "1100110001001" =>  data <= "11111111";  -- 1989 = FF
      when "1100110001010" =>  data <= "11111111";  -- 198A = FF
      when "1100110001011" =>  data <= "11111111";  -- 198B = FF
      when "1100110001100" =>  data <= "11111111";  -- 198C = FF
      when "1100110001101" =>  data <= "11111111";  -- 198D = FF
      when "1100110001110" =>  data <= "11111111";  -- 198E = FF
      when "1100110001111" =>  data <= "11111111";  -- 198F = FF
      when "1100110010000" =>  data <= "11111111";  -- 1990 = FF
      when "1100110010001" =>  data <= "11111111";  -- 1991 = FF
      when "1100110010010" =>  data <= "11111111";  -- 1992 = FF
      when "1100110010011" =>  data <= "11111111";  -- 1993 = FF
      when "1100110010100" =>  data <= "11111111";  -- 1994 = FF
      when "1100110010101" =>  data <= "11111111";  -- 1995 = FF
      when "1100110010110" =>  data <= "11111111";  -- 1996 = FF
      when "1100110010111" =>  data <= "11111111";  -- 1997 = FF
      when "1100110011000" =>  data <= "11111111";  -- 1998 = FF
      when "1100110011001" =>  data <= "11111111";  -- 1999 = FF
      when "1100110011010" =>  data <= "11111111";  -- 199A = FF
      when "1100110011011" =>  data <= "11111111";  -- 199B = FF
      when "1100110011100" =>  data <= "11111111";  -- 199C = FF
      when "1100110011101" =>  data <= "11111111";  -- 199D = FF
      when "1100110011110" =>  data <= "11111111";  -- 199E = FF
      when "1100110011111" =>  data <= "11111111";  -- 199F = FF
      when "1100110100000" =>  data <= "11111111";  -- 19A0 = FF
      when "1100110100001" =>  data <= "11111111";  -- 19A1 = FF
      when "1100110100010" =>  data <= "11111111";  -- 19A2 = FF
      when "1100110100011" =>  data <= "11111111";  -- 19A3 = FF
      when "1100110100100" =>  data <= "11111111";  -- 19A4 = FF
      when "1100110100101" =>  data <= "11111111";  -- 19A5 = FF
      when "1100110100110" =>  data <= "11111111";  -- 19A6 = FF
      when "1100110100111" =>  data <= "11111111";  -- 19A7 = FF
      when "1100110101000" =>  data <= "11111111";  -- 19A8 = FF
      when "1100110101001" =>  data <= "11111111";  -- 19A9 = FF
      when "1100110101010" =>  data <= "11111111";  -- 19AA = FF
      when "1100110101011" =>  data <= "11111111";  -- 19AB = FF
      when "1100110101100" =>  data <= "11111111";  -- 19AC = FF
      when "1100110101101" =>  data <= "11111111";  -- 19AD = FF
      when "1100110101110" =>  data <= "11111111";  -- 19AE = FF
      when "1100110101111" =>  data <= "11111111";  -- 19AF = FF
      when "1100110110000" =>  data <= "11111111";  -- 19B0 = FF
      when "1100110110001" =>  data <= "11111111";  -- 19B1 = FF
      when "1100110110010" =>  data <= "11111111";  -- 19B2 = FF
      when "1100110110011" =>  data <= "11111111";  -- 19B3 = FF
      when "1100110110100" =>  data <= "11111111";  -- 19B4 = FF
      when "1100110110101" =>  data <= "11111111";  -- 19B5 = FF
      when "1100110110110" =>  data <= "11111111";  -- 19B6 = FF
      when "1100110110111" =>  data <= "11111111";  -- 19B7 = FF
      when "1100110111000" =>  data <= "11111111";  -- 19B8 = FF
      when "1100110111001" =>  data <= "11111111";  -- 19B9 = FF
      when "1100110111010" =>  data <= "11111111";  -- 19BA = FF
      when "1100110111011" =>  data <= "11111111";  -- 19BB = FF
      when "1100110111100" =>  data <= "11111111";  -- 19BC = FF
      when "1100110111101" =>  data <= "11111111";  -- 19BD = FF
      when "1100110111110" =>  data <= "11111111";  -- 19BE = FF
      when "1100110111111" =>  data <= "11111111";  -- 19BF = FF
      when "1100111000000" =>  data <= "11111111";  -- 19C0 = FF
      when "1100111000001" =>  data <= "11111111";  -- 19C1 = FF
      when "1100111000010" =>  data <= "11111111";  -- 19C2 = FF
      when "1100111000011" =>  data <= "11111111";  -- 19C3 = FF
      when "1100111000100" =>  data <= "11111111";  -- 19C4 = FF
      when "1100111000101" =>  data <= "11111111";  -- 19C5 = FF
      when "1100111000110" =>  data <= "11111111";  -- 19C6 = FF
      when "1100111000111" =>  data <= "11111111";  -- 19C7 = FF
      when "1100111001000" =>  data <= "11111111";  -- 19C8 = FF
      when "1100111001001" =>  data <= "11111111";  -- 19C9 = FF
      when "1100111001010" =>  data <= "11111111";  -- 19CA = FF
      when "1100111001011" =>  data <= "11111111";  -- 19CB = FF
      when "1100111001100" =>  data <= "11111111";  -- 19CC = FF
      when "1100111001101" =>  data <= "11111111";  -- 19CD = FF
      when "1100111001110" =>  data <= "11111111";  -- 19CE = FF
      when "1100111001111" =>  data <= "11111111";  -- 19CF = FF
      when "1100111010000" =>  data <= "11111111";  -- 19D0 = FF
      when "1100111010001" =>  data <= "11111111";  -- 19D1 = FF
      when "1100111010010" =>  data <= "11111111";  -- 19D2 = FF
      when "1100111010011" =>  data <= "11111111";  -- 19D3 = FF
      when "1100111010100" =>  data <= "11111111";  -- 19D4 = FF
      when "1100111010101" =>  data <= "11111111";  -- 19D5 = FF
      when "1100111010110" =>  data <= "11111111";  -- 19D6 = FF
      when "1100111010111" =>  data <= "11111111";  -- 19D7 = FF
      when "1100111011000" =>  data <= "11111111";  -- 19D8 = FF
      when "1100111011001" =>  data <= "11111111";  -- 19D9 = FF
      when "1100111011010" =>  data <= "11111111";  -- 19DA = FF
      when "1100111011011" =>  data <= "11111111";  -- 19DB = FF
      when "1100111011100" =>  data <= "11111111";  -- 19DC = FF
      when "1100111011101" =>  data <= "11111111";  -- 19DD = FF
      when "1100111011110" =>  data <= "11111111";  -- 19DE = FF
      when "1100111011111" =>  data <= "11111111";  -- 19DF = FF
      when "1100111100000" =>  data <= "11111111";  -- 19E0 = FF
      when "1100111100001" =>  data <= "11111111";  -- 19E1 = FF
      when "1100111100010" =>  data <= "11111111";  -- 19E2 = FF
      when "1100111100011" =>  data <= "11111111";  -- 19E3 = FF
      when "1100111100100" =>  data <= "11111111";  -- 19E4 = FF
      when "1100111100101" =>  data <= "11111111";  -- 19E5 = FF
      when "1100111100110" =>  data <= "11111111";  -- 19E6 = FF
      when "1100111100111" =>  data <= "11111111";  -- 19E7 = FF
      when "1100111101000" =>  data <= "11111111";  -- 19E8 = FF
      when "1100111101001" =>  data <= "11111111";  -- 19E9 = FF
      when "1100111101010" =>  data <= "11111111";  -- 19EA = FF
      when "1100111101011" =>  data <= "11111111";  -- 19EB = FF
      when "1100111101100" =>  data <= "11111111";  -- 19EC = FF
      when "1100111101101" =>  data <= "11111111";  -- 19ED = FF
      when "1100111101110" =>  data <= "11111111";  -- 19EE = FF
      when "1100111101111" =>  data <= "11111111";  -- 19EF = FF
      when "1100111110000" =>  data <= "11111111";  -- 19F0 = FF
      when "1100111110001" =>  data <= "11111111";  -- 19F1 = FF
      when "1100111110010" =>  data <= "11111111";  -- 19F2 = FF
      when "1100111110011" =>  data <= "11111111";  -- 19F3 = FF
      when "1100111110100" =>  data <= "11111111";  -- 19F4 = FF
      when "1100111110101" =>  data <= "11111111";  -- 19F5 = FF
      when "1100111110110" =>  data <= "11111111";  -- 19F6 = FF
      when "1100111110111" =>  data <= "11111111";  -- 19F7 = FF
      when "1100111111000" =>  data <= "11111111";  -- 19F8 = FF
      when "1100111111001" =>  data <= "11111111";  -- 19F9 = FF
      when "1100111111010" =>  data <= "11111111";  -- 19FA = FF
      when "1100111111011" =>  data <= "11111111";  -- 19FB = FF
      when "1100111111100" =>  data <= "11111111";  -- 19FC = FF
      when "1100111111101" =>  data <= "11111111";  -- 19FD = FF
      when "1100111111110" =>  data <= "11111111";  -- 19FE = FF
      when "1100111111111" =>  data <= "11111111";  -- 19FF = FF
      when "1101000000000" =>  data <= "11111111";  -- 1A00 = FF
      when "1101000000001" =>  data <= "11111111";  -- 1A01 = FF
      when "1101000000010" =>  data <= "11111111";  -- 1A02 = FF
      when "1101000000011" =>  data <= "11111111";  -- 1A03 = FF
      when "1101000000100" =>  data <= "11111111";  -- 1A04 = FF
      when "1101000000101" =>  data <= "11111111";  -- 1A05 = FF
      when "1101000000110" =>  data <= "11111111";  -- 1A06 = FF
      when "1101000000111" =>  data <= "11111111";  -- 1A07 = FF
      when "1101000001000" =>  data <= "11111111";  -- 1A08 = FF
      when "1101000001001" =>  data <= "11111111";  -- 1A09 = FF
      when "1101000001010" =>  data <= "11111111";  -- 1A0A = FF
      when "1101000001011" =>  data <= "11111111";  -- 1A0B = FF
      when "1101000001100" =>  data <= "11111111";  -- 1A0C = FF
      when "1101000001101" =>  data <= "11111111";  -- 1A0D = FF
      when "1101000001110" =>  data <= "11111111";  -- 1A0E = FF
      when "1101000001111" =>  data <= "11111111";  -- 1A0F = FF
      when "1101000010000" =>  data <= "11111111";  -- 1A10 = FF
      when "1101000010001" =>  data <= "11111111";  -- 1A11 = FF
      when "1101000010010" =>  data <= "11111111";  -- 1A12 = FF
      when "1101000010011" =>  data <= "11111111";  -- 1A13 = FF
      when "1101000010100" =>  data <= "11111111";  -- 1A14 = FF
      when "1101000010101" =>  data <= "11111111";  -- 1A15 = FF
      when "1101000010110" =>  data <= "11111111";  -- 1A16 = FF
      when "1101000010111" =>  data <= "11111111";  -- 1A17 = FF
      when "1101000011000" =>  data <= "11111111";  -- 1A18 = FF
      when "1101000011001" =>  data <= "11111111";  -- 1A19 = FF
      when "1101000011010" =>  data <= "11111111";  -- 1A1A = FF
      when "1101000011011" =>  data <= "11111111";  -- 1A1B = FF
      when "1101000011100" =>  data <= "11111111";  -- 1A1C = FF
      when "1101000011101" =>  data <= "11111111";  -- 1A1D = FF
      when "1101000011110" =>  data <= "11111111";  -- 1A1E = FF
      when "1101000011111" =>  data <= "11111111";  -- 1A1F = FF
      when "1101000100000" =>  data <= "11111111";  -- 1A20 = FF
      when "1101000100001" =>  data <= "11111111";  -- 1A21 = FF
      when "1101000100010" =>  data <= "11111111";  -- 1A22 = FF
      when "1101000100011" =>  data <= "11111111";  -- 1A23 = FF
      when "1101000100100" =>  data <= "11111111";  -- 1A24 = FF
      when "1101000100101" =>  data <= "11111111";  -- 1A25 = FF
      when "1101000100110" =>  data <= "11111111";  -- 1A26 = FF
      when "1101000100111" =>  data <= "11111111";  -- 1A27 = FF
      when "1101000101000" =>  data <= "11111111";  -- 1A28 = FF
      when "1101000101001" =>  data <= "11111111";  -- 1A29 = FF
      when "1101000101010" =>  data <= "11111111";  -- 1A2A = FF
      when "1101000101011" =>  data <= "11111111";  -- 1A2B = FF
      when "1101000101100" =>  data <= "11111111";  -- 1A2C = FF
      when "1101000101101" =>  data <= "11111111";  -- 1A2D = FF
      when "1101000101110" =>  data <= "11111111";  -- 1A2E = FF
      when "1101000101111" =>  data <= "11111111";  -- 1A2F = FF
      when "1101000110000" =>  data <= "11111111";  -- 1A30 = FF
      when "1101000110001" =>  data <= "11111111";  -- 1A31 = FF
      when "1101000110010" =>  data <= "11111111";  -- 1A32 = FF
      when "1101000110011" =>  data <= "11111111";  -- 1A33 = FF
      when "1101000110100" =>  data <= "11111111";  -- 1A34 = FF
      when "1101000110101" =>  data <= "11111111";  -- 1A35 = FF
      when "1101000110110" =>  data <= "11111111";  -- 1A36 = FF
      when "1101000110111" =>  data <= "11111111";  -- 1A37 = FF
      when "1101000111000" =>  data <= "11111111";  -- 1A38 = FF
      when "1101000111001" =>  data <= "11111111";  -- 1A39 = FF
      when "1101000111010" =>  data <= "11111111";  -- 1A3A = FF
      when "1101000111011" =>  data <= "11111111";  -- 1A3B = FF
      when "1101000111100" =>  data <= "11111111";  -- 1A3C = FF
      when "1101000111101" =>  data <= "11111111";  -- 1A3D = FF
      when "1101000111110" =>  data <= "11111111";  -- 1A3E = FF
      when "1101000111111" =>  data <= "11111111";  -- 1A3F = FF
      when "1101001000000" =>  data <= "11111111";  -- 1A40 = FF
      when "1101001000001" =>  data <= "11111111";  -- 1A41 = FF
      when "1101001000010" =>  data <= "11111111";  -- 1A42 = FF
      when "1101001000011" =>  data <= "11111111";  -- 1A43 = FF
      when "1101001000100" =>  data <= "11111111";  -- 1A44 = FF
      when "1101001000101" =>  data <= "11111111";  -- 1A45 = FF
      when "1101001000110" =>  data <= "11111111";  -- 1A46 = FF
      when "1101001000111" =>  data <= "11111111";  -- 1A47 = FF
      when "1101001001000" =>  data <= "11111111";  -- 1A48 = FF
      when "1101001001001" =>  data <= "11111111";  -- 1A49 = FF
      when "1101001001010" =>  data <= "11111111";  -- 1A4A = FF
      when "1101001001011" =>  data <= "11111111";  -- 1A4B = FF
      when "1101001001100" =>  data <= "11111111";  -- 1A4C = FF
      when "1101001001101" =>  data <= "11111111";  -- 1A4D = FF
      when "1101001001110" =>  data <= "11111111";  -- 1A4E = FF
      when "1101001001111" =>  data <= "11111111";  -- 1A4F = FF
      when "1101001010000" =>  data <= "11111111";  -- 1A50 = FF
      when "1101001010001" =>  data <= "11111111";  -- 1A51 = FF
      when "1101001010010" =>  data <= "11111111";  -- 1A52 = FF
      when "1101001010011" =>  data <= "11111111";  -- 1A53 = FF
      when "1101001010100" =>  data <= "11111111";  -- 1A54 = FF
      when "1101001010101" =>  data <= "11111111";  -- 1A55 = FF
      when "1101001010110" =>  data <= "11111111";  -- 1A56 = FF
      when "1101001010111" =>  data <= "11111111";  -- 1A57 = FF
      when "1101001011000" =>  data <= "11111111";  -- 1A58 = FF
      when "1101001011001" =>  data <= "11111111";  -- 1A59 = FF
      when "1101001011010" =>  data <= "11111111";  -- 1A5A = FF
      when "1101001011011" =>  data <= "11111111";  -- 1A5B = FF
      when "1101001011100" =>  data <= "11111111";  -- 1A5C = FF
      when "1101001011101" =>  data <= "11111111";  -- 1A5D = FF
      when "1101001011110" =>  data <= "11111111";  -- 1A5E = FF
      when "1101001011111" =>  data <= "11111111";  -- 1A5F = FF
      when "1101001100000" =>  data <= "11111111";  -- 1A60 = FF
      when "1101001100001" =>  data <= "11111111";  -- 1A61 = FF
      when "1101001100010" =>  data <= "11111111";  -- 1A62 = FF
      when "1101001100011" =>  data <= "11111111";  -- 1A63 = FF
      when "1101001100100" =>  data <= "11111111";  -- 1A64 = FF
      when "1101001100101" =>  data <= "11111111";  -- 1A65 = FF
      when "1101001100110" =>  data <= "11111111";  -- 1A66 = FF
      when "1101001100111" =>  data <= "11111111";  -- 1A67 = FF
      when "1101001101000" =>  data <= "11111111";  -- 1A68 = FF
      when "1101001101001" =>  data <= "11111111";  -- 1A69 = FF
      when "1101001101010" =>  data <= "11111111";  -- 1A6A = FF
      when "1101001101011" =>  data <= "11111111";  -- 1A6B = FF
      when "1101001101100" =>  data <= "11111111";  -- 1A6C = FF
      when "1101001101101" =>  data <= "11111111";  -- 1A6D = FF
      when "1101001101110" =>  data <= "11111111";  -- 1A6E = FF
      when "1101001101111" =>  data <= "11111111";  -- 1A6F = FF
      when "1101001110000" =>  data <= "11111111";  -- 1A70 = FF
      when "1101001110001" =>  data <= "11111111";  -- 1A71 = FF
      when "1101001110010" =>  data <= "11111111";  -- 1A72 = FF
      when "1101001110011" =>  data <= "11111111";  -- 1A73 = FF
      when "1101001110100" =>  data <= "11111111";  -- 1A74 = FF
      when "1101001110101" =>  data <= "11111111";  -- 1A75 = FF
      when "1101001110110" =>  data <= "11111111";  -- 1A76 = FF
      when "1101001110111" =>  data <= "11111111";  -- 1A77 = FF
      when "1101001111000" =>  data <= "11111111";  -- 1A78 = FF
      when "1101001111001" =>  data <= "11111111";  -- 1A79 = FF
      when "1101001111010" =>  data <= "11111111";  -- 1A7A = FF
      when "1101001111011" =>  data <= "11111111";  -- 1A7B = FF
      when "1101001111100" =>  data <= "11111111";  -- 1A7C = FF
      when "1101001111101" =>  data <= "11111111";  -- 1A7D = FF
      when "1101001111110" =>  data <= "11111111";  -- 1A7E = FF
      when "1101001111111" =>  data <= "11111111";  -- 1A7F = FF
      when "1101010000000" =>  data <= "11111111";  -- 1A80 = FF
      when "1101010000001" =>  data <= "11111111";  -- 1A81 = FF
      when "1101010000010" =>  data <= "11111111";  -- 1A82 = FF
      when "1101010000011" =>  data <= "11111111";  -- 1A83 = FF
      when "1101010000100" =>  data <= "11111111";  -- 1A84 = FF
      when "1101010000101" =>  data <= "11111111";  -- 1A85 = FF
      when "1101010000110" =>  data <= "11111111";  -- 1A86 = FF
      when "1101010000111" =>  data <= "11111111";  -- 1A87 = FF
      when "1101010001000" =>  data <= "11111111";  -- 1A88 = FF
      when "1101010001001" =>  data <= "11111111";  -- 1A89 = FF
      when "1101010001010" =>  data <= "11111111";  -- 1A8A = FF
      when "1101010001011" =>  data <= "11111111";  -- 1A8B = FF
      when "1101010001100" =>  data <= "11111111";  -- 1A8C = FF
      when "1101010001101" =>  data <= "11111111";  -- 1A8D = FF
      when "1101010001110" =>  data <= "11111111";  -- 1A8E = FF
      when "1101010001111" =>  data <= "11111111";  -- 1A8F = FF
      when "1101010010000" =>  data <= "11111111";  -- 1A90 = FF
      when "1101010010001" =>  data <= "11111111";  -- 1A91 = FF
      when "1101010010010" =>  data <= "11111111";  -- 1A92 = FF
      when "1101010010011" =>  data <= "11111111";  -- 1A93 = FF
      when "1101010010100" =>  data <= "11111111";  -- 1A94 = FF
      when "1101010010101" =>  data <= "11111111";  -- 1A95 = FF
      when "1101010010110" =>  data <= "11111111";  -- 1A96 = FF
      when "1101010010111" =>  data <= "11111111";  -- 1A97 = FF
      when "1101010011000" =>  data <= "11111111";  -- 1A98 = FF
      when "1101010011001" =>  data <= "11111111";  -- 1A99 = FF
      when "1101010011010" =>  data <= "11111111";  -- 1A9A = FF
      when "1101010011011" =>  data <= "11111111";  -- 1A9B = FF
      when "1101010011100" =>  data <= "11111111";  -- 1A9C = FF
      when "1101010011101" =>  data <= "11111111";  -- 1A9D = FF
      when "1101010011110" =>  data <= "11111111";  -- 1A9E = FF
      when "1101010011111" =>  data <= "11111111";  -- 1A9F = FF
      when "1101010100000" =>  data <= "11111111";  -- 1AA0 = FF
      when "1101010100001" =>  data <= "11111111";  -- 1AA1 = FF
      when "1101010100010" =>  data <= "11111111";  -- 1AA2 = FF
      when "1101010100011" =>  data <= "11111111";  -- 1AA3 = FF
      when "1101010100100" =>  data <= "11111111";  -- 1AA4 = FF
      when "1101010100101" =>  data <= "11111111";  -- 1AA5 = FF
      when "1101010100110" =>  data <= "11111111";  -- 1AA6 = FF
      when "1101010100111" =>  data <= "11111111";  -- 1AA7 = FF
      when "1101010101000" =>  data <= "11111111";  -- 1AA8 = FF
      when "1101010101001" =>  data <= "11111111";  -- 1AA9 = FF
      when "1101010101010" =>  data <= "11111111";  -- 1AAA = FF
      when "1101010101011" =>  data <= "11111111";  -- 1AAB = FF
      when "1101010101100" =>  data <= "11111111";  -- 1AAC = FF
      when "1101010101101" =>  data <= "11111111";  -- 1AAD = FF
      when "1101010101110" =>  data <= "11111111";  -- 1AAE = FF
      when "1101010101111" =>  data <= "11111111";  -- 1AAF = FF
      when "1101010110000" =>  data <= "11111111";  -- 1AB0 = FF
      when "1101010110001" =>  data <= "11111111";  -- 1AB1 = FF
      when "1101010110010" =>  data <= "11111111";  -- 1AB2 = FF
      when "1101010110011" =>  data <= "11111111";  -- 1AB3 = FF
      when "1101010110100" =>  data <= "11111111";  -- 1AB4 = FF
      when "1101010110101" =>  data <= "11111111";  -- 1AB5 = FF
      when "1101010110110" =>  data <= "11111111";  -- 1AB6 = FF
      when "1101010110111" =>  data <= "11111111";  -- 1AB7 = FF
      when "1101010111000" =>  data <= "11111111";  -- 1AB8 = FF
      when "1101010111001" =>  data <= "11111111";  -- 1AB9 = FF
      when "1101010111010" =>  data <= "11111111";  -- 1ABA = FF
      when "1101010111011" =>  data <= "11111111";  -- 1ABB = FF
      when "1101010111100" =>  data <= "11111111";  -- 1ABC = FF
      when "1101010111101" =>  data <= "11111111";  -- 1ABD = FF
      when "1101010111110" =>  data <= "11111111";  -- 1ABE = FF
      when "1101010111111" =>  data <= "11111111";  -- 1ABF = FF
      when "1101011000000" =>  data <= "11111111";  -- 1AC0 = FF
      when "1101011000001" =>  data <= "11111111";  -- 1AC1 = FF
      when "1101011000010" =>  data <= "11111111";  -- 1AC2 = FF
      when "1101011000011" =>  data <= "11111111";  -- 1AC3 = FF
      when "1101011000100" =>  data <= "11111111";  -- 1AC4 = FF
      when "1101011000101" =>  data <= "11111111";  -- 1AC5 = FF
      when "1101011000110" =>  data <= "11111111";  -- 1AC6 = FF
      when "1101011000111" =>  data <= "11111111";  -- 1AC7 = FF
      when "1101011001000" =>  data <= "11111111";  -- 1AC8 = FF
      when "1101011001001" =>  data <= "11111111";  -- 1AC9 = FF
      when "1101011001010" =>  data <= "11111111";  -- 1ACA = FF
      when "1101011001011" =>  data <= "11111111";  -- 1ACB = FF
      when "1101011001100" =>  data <= "11111111";  -- 1ACC = FF
      when "1101011001101" =>  data <= "11111111";  -- 1ACD = FF
      when "1101011001110" =>  data <= "11111111";  -- 1ACE = FF
      when "1101011001111" =>  data <= "11111111";  -- 1ACF = FF
      when "1101011010000" =>  data <= "11111111";  -- 1AD0 = FF
      when "1101011010001" =>  data <= "11111111";  -- 1AD1 = FF
      when "1101011010010" =>  data <= "11111111";  -- 1AD2 = FF
      when "1101011010011" =>  data <= "11111111";  -- 1AD3 = FF
      when "1101011010100" =>  data <= "11111111";  -- 1AD4 = FF
      when "1101011010101" =>  data <= "11111111";  -- 1AD5 = FF
      when "1101011010110" =>  data <= "11111111";  -- 1AD6 = FF
      when "1101011010111" =>  data <= "11111111";  -- 1AD7 = FF
      when "1101011011000" =>  data <= "11111111";  -- 1AD8 = FF
      when "1101011011001" =>  data <= "11111111";  -- 1AD9 = FF
      when "1101011011010" =>  data <= "11111111";  -- 1ADA = FF
      when "1101011011011" =>  data <= "11111111";  -- 1ADB = FF
      when "1101011011100" =>  data <= "11111111";  -- 1ADC = FF
      when "1101011011101" =>  data <= "11111111";  -- 1ADD = FF
      when "1101011011110" =>  data <= "11111111";  -- 1ADE = FF
      when "1101011011111" =>  data <= "11111111";  -- 1ADF = FF
      when "1101011100000" =>  data <= "11111111";  -- 1AE0 = FF
      when "1101011100001" =>  data <= "11111111";  -- 1AE1 = FF
      when "1101011100010" =>  data <= "11111111";  -- 1AE2 = FF
      when "1101011100011" =>  data <= "11111111";  -- 1AE3 = FF
      when "1101011100100" =>  data <= "11111111";  -- 1AE4 = FF
      when "1101011100101" =>  data <= "11111111";  -- 1AE5 = FF
      when "1101011100110" =>  data <= "11111111";  -- 1AE6 = FF
      when "1101011100111" =>  data <= "11111111";  -- 1AE7 = FF
      when "1101011101000" =>  data <= "11111111";  -- 1AE8 = FF
      when "1101011101001" =>  data <= "11111111";  -- 1AE9 = FF
      when "1101011101010" =>  data <= "11111111";  -- 1AEA = FF
      when "1101011101011" =>  data <= "11111111";  -- 1AEB = FF
      when "1101011101100" =>  data <= "11111111";  -- 1AEC = FF
      when "1101011101101" =>  data <= "11111111";  -- 1AED = FF
      when "1101011101110" =>  data <= "11111111";  -- 1AEE = FF
      when "1101011101111" =>  data <= "11111111";  -- 1AEF = FF
      when "1101011110000" =>  data <= "11111111";  -- 1AF0 = FF
      when "1101011110001" =>  data <= "11111111";  -- 1AF1 = FF
      when "1101011110010" =>  data <= "11111111";  -- 1AF2 = FF
      when "1101011110011" =>  data <= "11111111";  -- 1AF3 = FF
      when "1101011110100" =>  data <= "11111111";  -- 1AF4 = FF
      when "1101011110101" =>  data <= "11111111";  -- 1AF5 = FF
      when "1101011110110" =>  data <= "11111111";  -- 1AF6 = FF
      when "1101011110111" =>  data <= "11111111";  -- 1AF7 = FF
      when "1101011111000" =>  data <= "11111111";  -- 1AF8 = FF
      when "1101011111001" =>  data <= "11111111";  -- 1AF9 = FF
      when "1101011111010" =>  data <= "11111111";  -- 1AFA = FF
      when "1101011111011" =>  data <= "11111111";  -- 1AFB = FF
      when "1101011111100" =>  data <= "11111111";  -- 1AFC = FF
      when "1101011111101" =>  data <= "11111111";  -- 1AFD = FF
      when "1101011111110" =>  data <= "11111111";  -- 1AFE = FF
      when "1101011111111" =>  data <= "11111111";  -- 1AFF = FF
      when "1101100000000" =>  data <= "11111111";  -- 1B00 = FF
      when "1101100000001" =>  data <= "11111111";  -- 1B01 = FF
      when "1101100000010" =>  data <= "11111111";  -- 1B02 = FF
      when "1101100000011" =>  data <= "11111111";  -- 1B03 = FF
      when "1101100000100" =>  data <= "11111111";  -- 1B04 = FF
      when "1101100000101" =>  data <= "11111111";  -- 1B05 = FF
      when "1101100000110" =>  data <= "11111111";  -- 1B06 = FF
      when "1101100000111" =>  data <= "11111111";  -- 1B07 = FF
      when "1101100001000" =>  data <= "11111111";  -- 1B08 = FF
      when "1101100001001" =>  data <= "11111111";  -- 1B09 = FF
      when "1101100001010" =>  data <= "11111111";  -- 1B0A = FF
      when "1101100001011" =>  data <= "11111111";  -- 1B0B = FF
      when "1101100001100" =>  data <= "11111111";  -- 1B0C = FF
      when "1101100001101" =>  data <= "11111111";  -- 1B0D = FF
      when "1101100001110" =>  data <= "11111111";  -- 1B0E = FF
      when "1101100001111" =>  data <= "11111111";  -- 1B0F = FF
      when "1101100010000" =>  data <= "11111111";  -- 1B10 = FF
      when "1101100010001" =>  data <= "11111111";  -- 1B11 = FF
      when "1101100010010" =>  data <= "11111111";  -- 1B12 = FF
      when "1101100010011" =>  data <= "11111111";  -- 1B13 = FF
      when "1101100010100" =>  data <= "11111111";  -- 1B14 = FF
      when "1101100010101" =>  data <= "11111111";  -- 1B15 = FF
      when "1101100010110" =>  data <= "11111111";  -- 1B16 = FF
      when "1101100010111" =>  data <= "11111111";  -- 1B17 = FF
      when "1101100011000" =>  data <= "11111111";  -- 1B18 = FF
      when "1101100011001" =>  data <= "11111111";  -- 1B19 = FF
      when "1101100011010" =>  data <= "11111111";  -- 1B1A = FF
      when "1101100011011" =>  data <= "11111111";  -- 1B1B = FF
      when "1101100011100" =>  data <= "11111111";  -- 1B1C = FF
      when "1101100011101" =>  data <= "11111111";  -- 1B1D = FF
      when "1101100011110" =>  data <= "11111111";  -- 1B1E = FF
      when "1101100011111" =>  data <= "11111111";  -- 1B1F = FF
      when "1101100100000" =>  data <= "11111111";  -- 1B20 = FF
      when "1101100100001" =>  data <= "11111111";  -- 1B21 = FF
      when "1101100100010" =>  data <= "11111111";  -- 1B22 = FF
      when "1101100100011" =>  data <= "11111111";  -- 1B23 = FF
      when "1101100100100" =>  data <= "11111111";  -- 1B24 = FF
      when "1101100100101" =>  data <= "11111111";  -- 1B25 = FF
      when "1101100100110" =>  data <= "11111111";  -- 1B26 = FF
      when "1101100100111" =>  data <= "11111111";  -- 1B27 = FF
      when "1101100101000" =>  data <= "11111111";  -- 1B28 = FF
      when "1101100101001" =>  data <= "11111111";  -- 1B29 = FF
      when "1101100101010" =>  data <= "11111111";  -- 1B2A = FF
      when "1101100101011" =>  data <= "11111111";  -- 1B2B = FF
      when "1101100101100" =>  data <= "11111111";  -- 1B2C = FF
      when "1101100101101" =>  data <= "11111111";  -- 1B2D = FF
      when "1101100101110" =>  data <= "11111111";  -- 1B2E = FF
      when "1101100101111" =>  data <= "11111111";  -- 1B2F = FF
      when "1101100110000" =>  data <= "11111111";  -- 1B30 = FF
      when "1101100110001" =>  data <= "11111111";  -- 1B31 = FF
      when "1101100110010" =>  data <= "11111111";  -- 1B32 = FF
      when "1101100110011" =>  data <= "11111111";  -- 1B33 = FF
      when "1101100110100" =>  data <= "11111111";  -- 1B34 = FF
      when "1101100110101" =>  data <= "11111111";  -- 1B35 = FF
      when "1101100110110" =>  data <= "11111111";  -- 1B36 = FF
      when "1101100110111" =>  data <= "11111111";  -- 1B37 = FF
      when "1101100111000" =>  data <= "11111111";  -- 1B38 = FF
      when "1101100111001" =>  data <= "11111111";  -- 1B39 = FF
      when "1101100111010" =>  data <= "11111111";  -- 1B3A = FF
      when "1101100111011" =>  data <= "11111111";  -- 1B3B = FF
      when "1101100111100" =>  data <= "11111111";  -- 1B3C = FF
      when "1101100111101" =>  data <= "11111111";  -- 1B3D = FF
      when "1101100111110" =>  data <= "11111111";  -- 1B3E = FF
      when "1101100111111" =>  data <= "11111111";  -- 1B3F = FF
      when "1101101000000" =>  data <= "11111111";  -- 1B40 = FF
      when "1101101000001" =>  data <= "11111111";  -- 1B41 = FF
      when "1101101000010" =>  data <= "11111111";  -- 1B42 = FF
      when "1101101000011" =>  data <= "11111111";  -- 1B43 = FF
      when "1101101000100" =>  data <= "11111111";  -- 1B44 = FF
      when "1101101000101" =>  data <= "11111111";  -- 1B45 = FF
      when "1101101000110" =>  data <= "11111111";  -- 1B46 = FF
      when "1101101000111" =>  data <= "11111111";  -- 1B47 = FF
      when "1101101001000" =>  data <= "11111111";  -- 1B48 = FF
      when "1101101001001" =>  data <= "11111111";  -- 1B49 = FF
      when "1101101001010" =>  data <= "11111111";  -- 1B4A = FF
      when "1101101001011" =>  data <= "11111111";  -- 1B4B = FF
      when "1101101001100" =>  data <= "11111111";  -- 1B4C = FF
      when "1101101001101" =>  data <= "11111111";  -- 1B4D = FF
      when "1101101001110" =>  data <= "11111111";  -- 1B4E = FF
      when "1101101001111" =>  data <= "11111111";  -- 1B4F = FF
      when "1101101010000" =>  data <= "11111111";  -- 1B50 = FF
      when "1101101010001" =>  data <= "11111111";  -- 1B51 = FF
      when "1101101010010" =>  data <= "11111111";  -- 1B52 = FF
      when "1101101010011" =>  data <= "11111111";  -- 1B53 = FF
      when "1101101010100" =>  data <= "11111111";  -- 1B54 = FF
      when "1101101010101" =>  data <= "11111111";  -- 1B55 = FF
      when "1101101010110" =>  data <= "11111111";  -- 1B56 = FF
      when "1101101010111" =>  data <= "11111111";  -- 1B57 = FF
      when "1101101011000" =>  data <= "11111111";  -- 1B58 = FF
      when "1101101011001" =>  data <= "11111111";  -- 1B59 = FF
      when "1101101011010" =>  data <= "11111111";  -- 1B5A = FF
      when "1101101011011" =>  data <= "11111111";  -- 1B5B = FF
      when "1101101011100" =>  data <= "11111111";  -- 1B5C = FF
      when "1101101011101" =>  data <= "11111111";  -- 1B5D = FF
      when "1101101011110" =>  data <= "11111111";  -- 1B5E = FF
      when "1101101011111" =>  data <= "11111111";  -- 1B5F = FF
      when "1101101100000" =>  data <= "11111111";  -- 1B60 = FF
      when "1101101100001" =>  data <= "11111111";  -- 1B61 = FF
      when "1101101100010" =>  data <= "11111111";  -- 1B62 = FF
      when "1101101100011" =>  data <= "11111111";  -- 1B63 = FF
      when "1101101100100" =>  data <= "11111111";  -- 1B64 = FF
      when "1101101100101" =>  data <= "11111111";  -- 1B65 = FF
      when "1101101100110" =>  data <= "11111111";  -- 1B66 = FF
      when "1101101100111" =>  data <= "11111111";  -- 1B67 = FF
      when "1101101101000" =>  data <= "11111111";  -- 1B68 = FF
      when "1101101101001" =>  data <= "11111111";  -- 1B69 = FF
      when "1101101101010" =>  data <= "11111111";  -- 1B6A = FF
      when "1101101101011" =>  data <= "11111111";  -- 1B6B = FF
      when "1101101101100" =>  data <= "11111111";  -- 1B6C = FF
      when "1101101101101" =>  data <= "11111111";  -- 1B6D = FF
      when "1101101101110" =>  data <= "11111111";  -- 1B6E = FF
      when "1101101101111" =>  data <= "11111111";  -- 1B6F = FF
      when "1101101110000" =>  data <= "11111111";  -- 1B70 = FF
      when "1101101110001" =>  data <= "11111111";  -- 1B71 = FF
      when "1101101110010" =>  data <= "11111111";  -- 1B72 = FF
      when "1101101110011" =>  data <= "11111111";  -- 1B73 = FF
      when "1101101110100" =>  data <= "11111111";  -- 1B74 = FF
      when "1101101110101" =>  data <= "11111111";  -- 1B75 = FF
      when "1101101110110" =>  data <= "11111111";  -- 1B76 = FF
      when "1101101110111" =>  data <= "11111111";  -- 1B77 = FF
      when "1101101111000" =>  data <= "11111111";  -- 1B78 = FF
      when "1101101111001" =>  data <= "11111111";  -- 1B79 = FF
      when "1101101111010" =>  data <= "11111111";  -- 1B7A = FF
      when "1101101111011" =>  data <= "11111111";  -- 1B7B = FF
      when "1101101111100" =>  data <= "11111111";  -- 1B7C = FF
      when "1101101111101" =>  data <= "11111111";  -- 1B7D = FF
      when "1101101111110" =>  data <= "11111111";  -- 1B7E = FF
      when "1101101111111" =>  data <= "11111111";  -- 1B7F = FF
      when "1101110000000" =>  data <= "11111111";  -- 1B80 = FF
      when "1101110000001" =>  data <= "11111111";  -- 1B81 = FF
      when "1101110000010" =>  data <= "11111111";  -- 1B82 = FF
      when "1101110000011" =>  data <= "11111111";  -- 1B83 = FF
      when "1101110000100" =>  data <= "11111111";  -- 1B84 = FF
      when "1101110000101" =>  data <= "11111111";  -- 1B85 = FF
      when "1101110000110" =>  data <= "11111111";  -- 1B86 = FF
      when "1101110000111" =>  data <= "11111111";  -- 1B87 = FF
      when "1101110001000" =>  data <= "11111111";  -- 1B88 = FF
      when "1101110001001" =>  data <= "11111111";  -- 1B89 = FF
      when "1101110001010" =>  data <= "11111111";  -- 1B8A = FF
      when "1101110001011" =>  data <= "11111111";  -- 1B8B = FF
      when "1101110001100" =>  data <= "11111111";  -- 1B8C = FF
      when "1101110001101" =>  data <= "11111111";  -- 1B8D = FF
      when "1101110001110" =>  data <= "11111111";  -- 1B8E = FF
      when "1101110001111" =>  data <= "11111111";  -- 1B8F = FF
      when "1101110010000" =>  data <= "11111111";  -- 1B90 = FF
      when "1101110010001" =>  data <= "11111111";  -- 1B91 = FF
      when "1101110010010" =>  data <= "11111111";  -- 1B92 = FF
      when "1101110010011" =>  data <= "11111111";  -- 1B93 = FF
      when "1101110010100" =>  data <= "11111111";  -- 1B94 = FF
      when "1101110010101" =>  data <= "11111111";  -- 1B95 = FF
      when "1101110010110" =>  data <= "11111111";  -- 1B96 = FF
      when "1101110010111" =>  data <= "11111111";  -- 1B97 = FF
      when "1101110011000" =>  data <= "11111111";  -- 1B98 = FF
      when "1101110011001" =>  data <= "11111111";  -- 1B99 = FF
      when "1101110011010" =>  data <= "11111111";  -- 1B9A = FF
      when "1101110011011" =>  data <= "11111111";  -- 1B9B = FF
      when "1101110011100" =>  data <= "11111111";  -- 1B9C = FF
      when "1101110011101" =>  data <= "11111111";  -- 1B9D = FF
      when "1101110011110" =>  data <= "11111111";  -- 1B9E = FF
      when "1101110011111" =>  data <= "11111111";  -- 1B9F = FF
      when "1101110100000" =>  data <= "11111111";  -- 1BA0 = FF
      when "1101110100001" =>  data <= "11111111";  -- 1BA1 = FF
      when "1101110100010" =>  data <= "11111111";  -- 1BA2 = FF
      when "1101110100011" =>  data <= "11111111";  -- 1BA3 = FF
      when "1101110100100" =>  data <= "11111111";  -- 1BA4 = FF
      when "1101110100101" =>  data <= "11111111";  -- 1BA5 = FF
      when "1101110100110" =>  data <= "11111111";  -- 1BA6 = FF
      when "1101110100111" =>  data <= "11111111";  -- 1BA7 = FF
      when "1101110101000" =>  data <= "11111111";  -- 1BA8 = FF
      when "1101110101001" =>  data <= "11111111";  -- 1BA9 = FF
      when "1101110101010" =>  data <= "11111111";  -- 1BAA = FF
      when "1101110101011" =>  data <= "11111111";  -- 1BAB = FF
      when "1101110101100" =>  data <= "11111111";  -- 1BAC = FF
      when "1101110101101" =>  data <= "11111111";  -- 1BAD = FF
      when "1101110101110" =>  data <= "11111111";  -- 1BAE = FF
      when "1101110101111" =>  data <= "11111111";  -- 1BAF = FF
      when "1101110110000" =>  data <= "11111111";  -- 1BB0 = FF
      when "1101110110001" =>  data <= "11111111";  -- 1BB1 = FF
      when "1101110110010" =>  data <= "11111111";  -- 1BB2 = FF
      when "1101110110011" =>  data <= "11111111";  -- 1BB3 = FF
      when "1101110110100" =>  data <= "11111111";  -- 1BB4 = FF
      when "1101110110101" =>  data <= "11111111";  -- 1BB5 = FF
      when "1101110110110" =>  data <= "11111111";  -- 1BB6 = FF
      when "1101110110111" =>  data <= "11111111";  -- 1BB7 = FF
      when "1101110111000" =>  data <= "11111111";  -- 1BB8 = FF
      when "1101110111001" =>  data <= "11111111";  -- 1BB9 = FF
      when "1101110111010" =>  data <= "11111111";  -- 1BBA = FF
      when "1101110111011" =>  data <= "11111111";  -- 1BBB = FF
      when "1101110111100" =>  data <= "11111111";  -- 1BBC = FF
      when "1101110111101" =>  data <= "11111111";  -- 1BBD = FF
      when "1101110111110" =>  data <= "11111111";  -- 1BBE = FF
      when "1101110111111" =>  data <= "11111111";  -- 1BBF = FF
      when "1101111000000" =>  data <= "11111111";  -- 1BC0 = FF
      when "1101111000001" =>  data <= "11111111";  -- 1BC1 = FF
      when "1101111000010" =>  data <= "11111111";  -- 1BC2 = FF
      when "1101111000011" =>  data <= "11111111";  -- 1BC3 = FF
      when "1101111000100" =>  data <= "11111111";  -- 1BC4 = FF
      when "1101111000101" =>  data <= "11111111";  -- 1BC5 = FF
      when "1101111000110" =>  data <= "11111111";  -- 1BC6 = FF
      when "1101111000111" =>  data <= "11111111";  -- 1BC7 = FF
      when "1101111001000" =>  data <= "11111111";  -- 1BC8 = FF
      when "1101111001001" =>  data <= "11111111";  -- 1BC9 = FF
      when "1101111001010" =>  data <= "11111111";  -- 1BCA = FF
      when "1101111001011" =>  data <= "11111111";  -- 1BCB = FF
      when "1101111001100" =>  data <= "11111111";  -- 1BCC = FF
      when "1101111001101" =>  data <= "11111111";  -- 1BCD = FF
      when "1101111001110" =>  data <= "11111111";  -- 1BCE = FF
      when "1101111001111" =>  data <= "11111111";  -- 1BCF = FF
      when "1101111010000" =>  data <= "11111111";  -- 1BD0 = FF
      when "1101111010001" =>  data <= "11111111";  -- 1BD1 = FF
      when "1101111010010" =>  data <= "11111111";  -- 1BD2 = FF
      when "1101111010011" =>  data <= "11111111";  -- 1BD3 = FF
      when "1101111010100" =>  data <= "11111111";  -- 1BD4 = FF
      when "1101111010101" =>  data <= "11111111";  -- 1BD5 = FF
      when "1101111010110" =>  data <= "11111111";  -- 1BD6 = FF
      when "1101111010111" =>  data <= "11111111";  -- 1BD7 = FF
      when "1101111011000" =>  data <= "11111111";  -- 1BD8 = FF
      when "1101111011001" =>  data <= "11111111";  -- 1BD9 = FF
      when "1101111011010" =>  data <= "11111111";  -- 1BDA = FF
      when "1101111011011" =>  data <= "11111111";  -- 1BDB = FF
      when "1101111011100" =>  data <= "11111111";  -- 1BDC = FF
      when "1101111011101" =>  data <= "11111111";  -- 1BDD = FF
      when "1101111011110" =>  data <= "11111111";  -- 1BDE = FF
      when "1101111011111" =>  data <= "11111111";  -- 1BDF = FF
      when "1101111100000" =>  data <= "11111111";  -- 1BE0 = FF
      when "1101111100001" =>  data <= "11111111";  -- 1BE1 = FF
      when "1101111100010" =>  data <= "11111111";  -- 1BE2 = FF
      when "1101111100011" =>  data <= "11111111";  -- 1BE3 = FF
      when "1101111100100" =>  data <= "11111111";  -- 1BE4 = FF
      when "1101111100101" =>  data <= "11111111";  -- 1BE5 = FF
      when "1101111100110" =>  data <= "11111111";  -- 1BE6 = FF
      when "1101111100111" =>  data <= "11111111";  -- 1BE7 = FF
      when "1101111101000" =>  data <= "11111111";  -- 1BE8 = FF
      when "1101111101001" =>  data <= "11111111";  -- 1BE9 = FF
      when "1101111101010" =>  data <= "11111111";  -- 1BEA = FF
      when "1101111101011" =>  data <= "11111111";  -- 1BEB = FF
      when "1101111101100" =>  data <= "11111111";  -- 1BEC = FF
      when "1101111101101" =>  data <= "11111111";  -- 1BED = FF
      when "1101111101110" =>  data <= "11111111";  -- 1BEE = FF
      when "1101111101111" =>  data <= "11111111";  -- 1BEF = FF
      when "1101111110000" =>  data <= "11111111";  -- 1BF0 = FF
      when "1101111110001" =>  data <= "11111111";  -- 1BF1 = FF
      when "1101111110010" =>  data <= "11111111";  -- 1BF2 = FF
      when "1101111110011" =>  data <= "11111111";  -- 1BF3 = FF
      when "1101111110100" =>  data <= "11111111";  -- 1BF4 = FF
      when "1101111110101" =>  data <= "11111111";  -- 1BF5 = FF
      when "1101111110110" =>  data <= "11111111";  -- 1BF6 = FF
      when "1101111110111" =>  data <= "11111111";  -- 1BF7 = FF
      when "1101111111000" =>  data <= "11111111";  -- 1BF8 = FF
      when "1101111111001" =>  data <= "11111111";  -- 1BF9 = FF
      when "1101111111010" =>  data <= "11111111";  -- 1BFA = FF
      when "1101111111011" =>  data <= "11111111";  -- 1BFB = FF
      when "1101111111100" =>  data <= "11111111";  -- 1BFC = FF
      when "1101111111101" =>  data <= "11111111";  -- 1BFD = FF
      when "1101111111110" =>  data <= "11111111";  -- 1BFE = FF
      when "1101111111111" =>  data <= "11111111";  -- 1BFF = FF
      when "1110000000000" =>  data <= "11111111";  -- 1C00 = FF
      when "1110000000001" =>  data <= "11111111";  -- 1C01 = FF
      when "1110000000010" =>  data <= "11111111";  -- 1C02 = FF
      when "1110000000011" =>  data <= "11111111";  -- 1C03 = FF
      when "1110000000100" =>  data <= "11111111";  -- 1C04 = FF
      when "1110000000101" =>  data <= "11111111";  -- 1C05 = FF
      when "1110000000110" =>  data <= "11111111";  -- 1C06 = FF
      when "1110000000111" =>  data <= "11111111";  -- 1C07 = FF
      when "1110000001000" =>  data <= "11111111";  -- 1C08 = FF
      when "1110000001001" =>  data <= "11111111";  -- 1C09 = FF
      when "1110000001010" =>  data <= "11111111";  -- 1C0A = FF
      when "1110000001011" =>  data <= "11111111";  -- 1C0B = FF
      when "1110000001100" =>  data <= "11111111";  -- 1C0C = FF
      when "1110000001101" =>  data <= "11111111";  -- 1C0D = FF
      when "1110000001110" =>  data <= "11111111";  -- 1C0E = FF
      when "1110000001111" =>  data <= "11111111";  -- 1C0F = FF
      when "1110000010000" =>  data <= "11111111";  -- 1C10 = FF
      when "1110000010001" =>  data <= "11111111";  -- 1C11 = FF
      when "1110000010010" =>  data <= "11111111";  -- 1C12 = FF
      when "1110000010011" =>  data <= "11111111";  -- 1C13 = FF
      when "1110000010100" =>  data <= "11111111";  -- 1C14 = FF
      when "1110000010101" =>  data <= "11111111";  -- 1C15 = FF
      when "1110000010110" =>  data <= "11111111";  -- 1C16 = FF
      when "1110000010111" =>  data <= "11111111";  -- 1C17 = FF
      when "1110000011000" =>  data <= "11111111";  -- 1C18 = FF
      when "1110000011001" =>  data <= "11111111";  -- 1C19 = FF
      when "1110000011010" =>  data <= "11111111";  -- 1C1A = FF
      when "1110000011011" =>  data <= "11111111";  -- 1C1B = FF
      when "1110000011100" =>  data <= "11111111";  -- 1C1C = FF
      when "1110000011101" =>  data <= "11111111";  -- 1C1D = FF
      when "1110000011110" =>  data <= "11111111";  -- 1C1E = FF
      when "1110000011111" =>  data <= "11111111";  -- 1C1F = FF
      when "1110000100000" =>  data <= "11111111";  -- 1C20 = FF
      when "1110000100001" =>  data <= "11111111";  -- 1C21 = FF
      when "1110000100010" =>  data <= "11111111";  -- 1C22 = FF
      when "1110000100011" =>  data <= "11111111";  -- 1C23 = FF
      when "1110000100100" =>  data <= "11111111";  -- 1C24 = FF
      when "1110000100101" =>  data <= "11111111";  -- 1C25 = FF
      when "1110000100110" =>  data <= "11111111";  -- 1C26 = FF
      when "1110000100111" =>  data <= "11111111";  -- 1C27 = FF
      when "1110000101000" =>  data <= "11111111";  -- 1C28 = FF
      when "1110000101001" =>  data <= "11111111";  -- 1C29 = FF
      when "1110000101010" =>  data <= "11111111";  -- 1C2A = FF
      when "1110000101011" =>  data <= "11111111";  -- 1C2B = FF
      when "1110000101100" =>  data <= "11111111";  -- 1C2C = FF
      when "1110000101101" =>  data <= "11111111";  -- 1C2D = FF
      when "1110000101110" =>  data <= "11111111";  -- 1C2E = FF
      when "1110000101111" =>  data <= "11111111";  -- 1C2F = FF
      when "1110000110000" =>  data <= "11111111";  -- 1C30 = FF
      when "1110000110001" =>  data <= "11111111";  -- 1C31 = FF
      when "1110000110010" =>  data <= "11111111";  -- 1C32 = FF
      when "1110000110011" =>  data <= "11111111";  -- 1C33 = FF
      when "1110000110100" =>  data <= "11111111";  -- 1C34 = FF
      when "1110000110101" =>  data <= "11111111";  -- 1C35 = FF
      when "1110000110110" =>  data <= "11111111";  -- 1C36 = FF
      when "1110000110111" =>  data <= "11111111";  -- 1C37 = FF
      when "1110000111000" =>  data <= "11111111";  -- 1C38 = FF
      when "1110000111001" =>  data <= "11111111";  -- 1C39 = FF
      when "1110000111010" =>  data <= "11111111";  -- 1C3A = FF
      when "1110000111011" =>  data <= "11111111";  -- 1C3B = FF
      when "1110000111100" =>  data <= "11111111";  -- 1C3C = FF
      when "1110000111101" =>  data <= "11111111";  -- 1C3D = FF
      when "1110000111110" =>  data <= "11111111";  -- 1C3E = FF
      when "1110000111111" =>  data <= "11111111";  -- 1C3F = FF
      when "1110001000000" =>  data <= "11111111";  -- 1C40 = FF
      when "1110001000001" =>  data <= "11111111";  -- 1C41 = FF
      when "1110001000010" =>  data <= "11111111";  -- 1C42 = FF
      when "1110001000011" =>  data <= "11111111";  -- 1C43 = FF
      when "1110001000100" =>  data <= "11111111";  -- 1C44 = FF
      when "1110001000101" =>  data <= "11111111";  -- 1C45 = FF
      when "1110001000110" =>  data <= "11111111";  -- 1C46 = FF
      when "1110001000111" =>  data <= "11111111";  -- 1C47 = FF
      when "1110001001000" =>  data <= "11111111";  -- 1C48 = FF
      when "1110001001001" =>  data <= "11111111";  -- 1C49 = FF
      when "1110001001010" =>  data <= "11111111";  -- 1C4A = FF
      when "1110001001011" =>  data <= "11111111";  -- 1C4B = FF
      when "1110001001100" =>  data <= "11111111";  -- 1C4C = FF
      when "1110001001101" =>  data <= "11111111";  -- 1C4D = FF
      when "1110001001110" =>  data <= "11111111";  -- 1C4E = FF
      when "1110001001111" =>  data <= "11111111";  -- 1C4F = FF
      when "1110001010000" =>  data <= "11111111";  -- 1C50 = FF
      when "1110001010001" =>  data <= "11111111";  -- 1C51 = FF
      when "1110001010010" =>  data <= "11111111";  -- 1C52 = FF
      when "1110001010011" =>  data <= "11111111";  -- 1C53 = FF
      when "1110001010100" =>  data <= "11111111";  -- 1C54 = FF
      when "1110001010101" =>  data <= "11111111";  -- 1C55 = FF
      when "1110001010110" =>  data <= "11111111";  -- 1C56 = FF
      when "1110001010111" =>  data <= "11111111";  -- 1C57 = FF
      when "1110001011000" =>  data <= "11111111";  -- 1C58 = FF
      when "1110001011001" =>  data <= "11111111";  -- 1C59 = FF
      when "1110001011010" =>  data <= "11111111";  -- 1C5A = FF
      when "1110001011011" =>  data <= "11111111";  -- 1C5B = FF
      when "1110001011100" =>  data <= "11111111";  -- 1C5C = FF
      when "1110001011101" =>  data <= "11111111";  -- 1C5D = FF
      when "1110001011110" =>  data <= "11111111";  -- 1C5E = FF
      when "1110001011111" =>  data <= "11111111";  -- 1C5F = FF
      when "1110001100000" =>  data <= "11111111";  -- 1C60 = FF
      when "1110001100001" =>  data <= "11111111";  -- 1C61 = FF
      when "1110001100010" =>  data <= "11111111";  -- 1C62 = FF
      when "1110001100011" =>  data <= "11111111";  -- 1C63 = FF
      when "1110001100100" =>  data <= "11111111";  -- 1C64 = FF
      when "1110001100101" =>  data <= "11111111";  -- 1C65 = FF
      when "1110001100110" =>  data <= "11111111";  -- 1C66 = FF
      when "1110001100111" =>  data <= "11111111";  -- 1C67 = FF
      when "1110001101000" =>  data <= "11111111";  -- 1C68 = FF
      when "1110001101001" =>  data <= "11111111";  -- 1C69 = FF
      when "1110001101010" =>  data <= "11111111";  -- 1C6A = FF
      when "1110001101011" =>  data <= "11111111";  -- 1C6B = FF
      when "1110001101100" =>  data <= "11111111";  -- 1C6C = FF
      when "1110001101101" =>  data <= "11111111";  -- 1C6D = FF
      when "1110001101110" =>  data <= "11111111";  -- 1C6E = FF
      when "1110001101111" =>  data <= "11111111";  -- 1C6F = FF
      when "1110001110000" =>  data <= "11111111";  -- 1C70 = FF
      when "1110001110001" =>  data <= "11111111";  -- 1C71 = FF
      when "1110001110010" =>  data <= "11111111";  -- 1C72 = FF
      when "1110001110011" =>  data <= "11111111";  -- 1C73 = FF
      when "1110001110100" =>  data <= "11111111";  -- 1C74 = FF
      when "1110001110101" =>  data <= "11111111";  -- 1C75 = FF
      when "1110001110110" =>  data <= "11111111";  -- 1C76 = FF
      when "1110001110111" =>  data <= "11111111";  -- 1C77 = FF
      when "1110001111000" =>  data <= "11111111";  -- 1C78 = FF
      when "1110001111001" =>  data <= "11111111";  -- 1C79 = FF
      when "1110001111010" =>  data <= "11111111";  -- 1C7A = FF
      when "1110001111011" =>  data <= "11111111";  -- 1C7B = FF
      when "1110001111100" =>  data <= "11111111";  -- 1C7C = FF
      when "1110001111101" =>  data <= "11111111";  -- 1C7D = FF
      when "1110001111110" =>  data <= "11111111";  -- 1C7E = FF
      when "1110001111111" =>  data <= "11111111";  -- 1C7F = FF
      when "1110010000000" =>  data <= "11111111";  -- 1C80 = FF
      when "1110010000001" =>  data <= "11111111";  -- 1C81 = FF
      when "1110010000010" =>  data <= "11111111";  -- 1C82 = FF
      when "1110010000011" =>  data <= "11111111";  -- 1C83 = FF
      when "1110010000100" =>  data <= "11111111";  -- 1C84 = FF
      when "1110010000101" =>  data <= "11111111";  -- 1C85 = FF
      when "1110010000110" =>  data <= "11111111";  -- 1C86 = FF
      when "1110010000111" =>  data <= "11111111";  -- 1C87 = FF
      when "1110010001000" =>  data <= "11111111";  -- 1C88 = FF
      when "1110010001001" =>  data <= "11111111";  -- 1C89 = FF
      when "1110010001010" =>  data <= "11111111";  -- 1C8A = FF
      when "1110010001011" =>  data <= "11111111";  -- 1C8B = FF
      when "1110010001100" =>  data <= "11111111";  -- 1C8C = FF
      when "1110010001101" =>  data <= "11111111";  -- 1C8D = FF
      when "1110010001110" =>  data <= "11111111";  -- 1C8E = FF
      when "1110010001111" =>  data <= "11111111";  -- 1C8F = FF
      when "1110010010000" =>  data <= "11111111";  -- 1C90 = FF
      when "1110010010001" =>  data <= "11111111";  -- 1C91 = FF
      when "1110010010010" =>  data <= "11111111";  -- 1C92 = FF
      when "1110010010011" =>  data <= "11111111";  -- 1C93 = FF
      when "1110010010100" =>  data <= "11111111";  -- 1C94 = FF
      when "1110010010101" =>  data <= "11111111";  -- 1C95 = FF
      when "1110010010110" =>  data <= "11111111";  -- 1C96 = FF
      when "1110010010111" =>  data <= "11111111";  -- 1C97 = FF
      when "1110010011000" =>  data <= "11111111";  -- 1C98 = FF
      when "1110010011001" =>  data <= "11111111";  -- 1C99 = FF
      when "1110010011010" =>  data <= "11111111";  -- 1C9A = FF
      when "1110010011011" =>  data <= "11111111";  -- 1C9B = FF
      when "1110010011100" =>  data <= "11111111";  -- 1C9C = FF
      when "1110010011101" =>  data <= "11111111";  -- 1C9D = FF
      when "1110010011110" =>  data <= "11111111";  -- 1C9E = FF
      when "1110010011111" =>  data <= "11111111";  -- 1C9F = FF
      when "1110010100000" =>  data <= "11111111";  -- 1CA0 = FF
      when "1110010100001" =>  data <= "11111111";  -- 1CA1 = FF
      when "1110010100010" =>  data <= "11111111";  -- 1CA2 = FF
      when "1110010100011" =>  data <= "11111111";  -- 1CA3 = FF
      when "1110010100100" =>  data <= "11111111";  -- 1CA4 = FF
      when "1110010100101" =>  data <= "11111111";  -- 1CA5 = FF
      when "1110010100110" =>  data <= "11111111";  -- 1CA6 = FF
      when "1110010100111" =>  data <= "11111111";  -- 1CA7 = FF
      when "1110010101000" =>  data <= "11111111";  -- 1CA8 = FF
      when "1110010101001" =>  data <= "11111111";  -- 1CA9 = FF
      when "1110010101010" =>  data <= "11111111";  -- 1CAA = FF
      when "1110010101011" =>  data <= "11111111";  -- 1CAB = FF
      when "1110010101100" =>  data <= "11111111";  -- 1CAC = FF
      when "1110010101101" =>  data <= "11111111";  -- 1CAD = FF
      when "1110010101110" =>  data <= "11111111";  -- 1CAE = FF
      when "1110010101111" =>  data <= "11111111";  -- 1CAF = FF
      when "1110010110000" =>  data <= "11111111";  -- 1CB0 = FF
      when "1110010110001" =>  data <= "11111111";  -- 1CB1 = FF
      when "1110010110010" =>  data <= "11111111";  -- 1CB2 = FF
      when "1110010110011" =>  data <= "11111111";  -- 1CB3 = FF
      when "1110010110100" =>  data <= "11111111";  -- 1CB4 = FF
      when "1110010110101" =>  data <= "11111111";  -- 1CB5 = FF
      when "1110010110110" =>  data <= "11111111";  -- 1CB6 = FF
      when "1110010110111" =>  data <= "11111111";  -- 1CB7 = FF
      when "1110010111000" =>  data <= "11111111";  -- 1CB8 = FF
      when "1110010111001" =>  data <= "11111111";  -- 1CB9 = FF
      when "1110010111010" =>  data <= "11111111";  -- 1CBA = FF
      when "1110010111011" =>  data <= "11111111";  -- 1CBB = FF
      when "1110010111100" =>  data <= "11111111";  -- 1CBC = FF
      when "1110010111101" =>  data <= "11111111";  -- 1CBD = FF
      when "1110010111110" =>  data <= "11111111";  -- 1CBE = FF
      when "1110010111111" =>  data <= "11111111";  -- 1CBF = FF
      when "1110011000000" =>  data <= "11111111";  -- 1CC0 = FF
      when "1110011000001" =>  data <= "11111111";  -- 1CC1 = FF
      when "1110011000010" =>  data <= "11111111";  -- 1CC2 = FF
      when "1110011000011" =>  data <= "11111111";  -- 1CC3 = FF
      when "1110011000100" =>  data <= "11111111";  -- 1CC4 = FF
      when "1110011000101" =>  data <= "11111111";  -- 1CC5 = FF
      when "1110011000110" =>  data <= "11111111";  -- 1CC6 = FF
      when "1110011000111" =>  data <= "11111111";  -- 1CC7 = FF
      when "1110011001000" =>  data <= "11111111";  -- 1CC8 = FF
      when "1110011001001" =>  data <= "11111111";  -- 1CC9 = FF
      when "1110011001010" =>  data <= "11111111";  -- 1CCA = FF
      when "1110011001011" =>  data <= "11111111";  -- 1CCB = FF
      when "1110011001100" =>  data <= "11111111";  -- 1CCC = FF
      when "1110011001101" =>  data <= "11111111";  -- 1CCD = FF
      when "1110011001110" =>  data <= "11111111";  -- 1CCE = FF
      when "1110011001111" =>  data <= "11111111";  -- 1CCF = FF
      when "1110011010000" =>  data <= "11111111";  -- 1CD0 = FF
      when "1110011010001" =>  data <= "11111111";  -- 1CD1 = FF
      when "1110011010010" =>  data <= "11111111";  -- 1CD2 = FF
      when "1110011010011" =>  data <= "11111111";  -- 1CD3 = FF
      when "1110011010100" =>  data <= "11111111";  -- 1CD4 = FF
      when "1110011010101" =>  data <= "11111111";  -- 1CD5 = FF
      when "1110011010110" =>  data <= "11111111";  -- 1CD6 = FF
      when "1110011010111" =>  data <= "11111111";  -- 1CD7 = FF
      when "1110011011000" =>  data <= "11111111";  -- 1CD8 = FF
      when "1110011011001" =>  data <= "11111111";  -- 1CD9 = FF
      when "1110011011010" =>  data <= "11111111";  -- 1CDA = FF
      when "1110011011011" =>  data <= "11111111";  -- 1CDB = FF
      when "1110011011100" =>  data <= "11111111";  -- 1CDC = FF
      when "1110011011101" =>  data <= "11111111";  -- 1CDD = FF
      when "1110011011110" =>  data <= "11111111";  -- 1CDE = FF
      when "1110011011111" =>  data <= "11111111";  -- 1CDF = FF
      when "1110011100000" =>  data <= "11111111";  -- 1CE0 = FF
      when "1110011100001" =>  data <= "11111111";  -- 1CE1 = FF
      when "1110011100010" =>  data <= "11111111";  -- 1CE2 = FF
      when "1110011100011" =>  data <= "11111111";  -- 1CE3 = FF
      when "1110011100100" =>  data <= "11111111";  -- 1CE4 = FF
      when "1110011100101" =>  data <= "11111111";  -- 1CE5 = FF
      when "1110011100110" =>  data <= "11111111";  -- 1CE6 = FF
      when "1110011100111" =>  data <= "11111111";  -- 1CE7 = FF
      when "1110011101000" =>  data <= "11111111";  -- 1CE8 = FF
      when "1110011101001" =>  data <= "11111111";  -- 1CE9 = FF
      when "1110011101010" =>  data <= "11111111";  -- 1CEA = FF
      when "1110011101011" =>  data <= "11111111";  -- 1CEB = FF
      when "1110011101100" =>  data <= "11111111";  -- 1CEC = FF
      when "1110011101101" =>  data <= "11111111";  -- 1CED = FF
      when "1110011101110" =>  data <= "11111111";  -- 1CEE = FF
      when "1110011101111" =>  data <= "11111111";  -- 1CEF = FF
      when "1110011110000" =>  data <= "11111111";  -- 1CF0 = FF
      when "1110011110001" =>  data <= "11111111";  -- 1CF1 = FF
      when "1110011110010" =>  data <= "11111111";  -- 1CF2 = FF
      when "1110011110011" =>  data <= "11111111";  -- 1CF3 = FF
      when "1110011110100" =>  data <= "11111111";  -- 1CF4 = FF
      when "1110011110101" =>  data <= "11111111";  -- 1CF5 = FF
      when "1110011110110" =>  data <= "11111111";  -- 1CF6 = FF
      when "1110011110111" =>  data <= "11111111";  -- 1CF7 = FF
      when "1110011111000" =>  data <= "11111111";  -- 1CF8 = FF
      when "1110011111001" =>  data <= "11111111";  -- 1CF9 = FF
      when "1110011111010" =>  data <= "11111111";  -- 1CFA = FF
      when "1110011111011" =>  data <= "11111111";  -- 1CFB = FF
      when "1110011111100" =>  data <= "11111111";  -- 1CFC = FF
      when "1110011111101" =>  data <= "11111111";  -- 1CFD = FF
      when "1110011111110" =>  data <= "11111111";  -- 1CFE = FF
      when "1110011111111" =>  data <= "11111111";  -- 1CFF = FF
      when "1110100000000" =>  data <= "11111111";  -- 1D00 = FF
      when "1110100000001" =>  data <= "11111111";  -- 1D01 = FF
      when "1110100000010" =>  data <= "11111111";  -- 1D02 = FF
      when "1110100000011" =>  data <= "11111111";  -- 1D03 = FF
      when "1110100000100" =>  data <= "11111111";  -- 1D04 = FF
      when "1110100000101" =>  data <= "11111111";  -- 1D05 = FF
      when "1110100000110" =>  data <= "11111111";  -- 1D06 = FF
      when "1110100000111" =>  data <= "11111111";  -- 1D07 = FF
      when "1110100001000" =>  data <= "11111111";  -- 1D08 = FF
      when "1110100001001" =>  data <= "11111111";  -- 1D09 = FF
      when "1110100001010" =>  data <= "11111111";  -- 1D0A = FF
      when "1110100001011" =>  data <= "11111111";  -- 1D0B = FF
      when "1110100001100" =>  data <= "11111111";  -- 1D0C = FF
      when "1110100001101" =>  data <= "11111111";  -- 1D0D = FF
      when "1110100001110" =>  data <= "11111111";  -- 1D0E = FF
      when "1110100001111" =>  data <= "11111111";  -- 1D0F = FF
      when "1110100010000" =>  data <= "11111111";  -- 1D10 = FF
      when "1110100010001" =>  data <= "11111111";  -- 1D11 = FF
      when "1110100010010" =>  data <= "11111111";  -- 1D12 = FF
      when "1110100010011" =>  data <= "11111111";  -- 1D13 = FF
      when "1110100010100" =>  data <= "11111111";  -- 1D14 = FF
      when "1110100010101" =>  data <= "11111111";  -- 1D15 = FF
      when "1110100010110" =>  data <= "11111111";  -- 1D16 = FF
      when "1110100010111" =>  data <= "11111111";  -- 1D17 = FF
      when "1110100011000" =>  data <= "11111111";  -- 1D18 = FF
      when "1110100011001" =>  data <= "11111111";  -- 1D19 = FF
      when "1110100011010" =>  data <= "11111111";  -- 1D1A = FF
      when "1110100011011" =>  data <= "11111111";  -- 1D1B = FF
      when "1110100011100" =>  data <= "11111111";  -- 1D1C = FF
      when "1110100011101" =>  data <= "11111111";  -- 1D1D = FF
      when "1110100011110" =>  data <= "11111111";  -- 1D1E = FF
      when "1110100011111" =>  data <= "11111111";  -- 1D1F = FF
      when "1110100100000" =>  data <= "11111111";  -- 1D20 = FF
      when "1110100100001" =>  data <= "11111111";  -- 1D21 = FF
      when "1110100100010" =>  data <= "11111111";  -- 1D22 = FF
      when "1110100100011" =>  data <= "11111111";  -- 1D23 = FF
      when "1110100100100" =>  data <= "11111111";  -- 1D24 = FF
      when "1110100100101" =>  data <= "11111111";  -- 1D25 = FF
      when "1110100100110" =>  data <= "11111111";  -- 1D26 = FF
      when "1110100100111" =>  data <= "11111111";  -- 1D27 = FF
      when "1110100101000" =>  data <= "11111111";  -- 1D28 = FF
      when "1110100101001" =>  data <= "11111111";  -- 1D29 = FF
      when "1110100101010" =>  data <= "11111111";  -- 1D2A = FF
      when "1110100101011" =>  data <= "11111111";  -- 1D2B = FF
      when "1110100101100" =>  data <= "11111111";  -- 1D2C = FF
      when "1110100101101" =>  data <= "11111111";  -- 1D2D = FF
      when "1110100101110" =>  data <= "11111111";  -- 1D2E = FF
      when "1110100101111" =>  data <= "11111111";  -- 1D2F = FF
      when "1110100110000" =>  data <= "11111111";  -- 1D30 = FF
      when "1110100110001" =>  data <= "11111111";  -- 1D31 = FF
      when "1110100110010" =>  data <= "11111111";  -- 1D32 = FF
      when "1110100110011" =>  data <= "11111111";  -- 1D33 = FF
      when "1110100110100" =>  data <= "11111111";  -- 1D34 = FF
      when "1110100110101" =>  data <= "11111111";  -- 1D35 = FF
      when "1110100110110" =>  data <= "11111111";  -- 1D36 = FF
      when "1110100110111" =>  data <= "11111111";  -- 1D37 = FF
      when "1110100111000" =>  data <= "11111111";  -- 1D38 = FF
      when "1110100111001" =>  data <= "11111111";  -- 1D39 = FF
      when "1110100111010" =>  data <= "11111111";  -- 1D3A = FF
      when "1110100111011" =>  data <= "11111111";  -- 1D3B = FF
      when "1110100111100" =>  data <= "11111111";  -- 1D3C = FF
      when "1110100111101" =>  data <= "11111111";  -- 1D3D = FF
      when "1110100111110" =>  data <= "11111111";  -- 1D3E = FF
      when "1110100111111" =>  data <= "11111111";  -- 1D3F = FF
      when "1110101000000" =>  data <= "11111111";  -- 1D40 = FF
      when "1110101000001" =>  data <= "11111111";  -- 1D41 = FF
      when "1110101000010" =>  data <= "11111111";  -- 1D42 = FF
      when "1110101000011" =>  data <= "11111111";  -- 1D43 = FF
      when "1110101000100" =>  data <= "11111111";  -- 1D44 = FF
      when "1110101000101" =>  data <= "11111111";  -- 1D45 = FF
      when "1110101000110" =>  data <= "11111111";  -- 1D46 = FF
      when "1110101000111" =>  data <= "11111111";  -- 1D47 = FF
      when "1110101001000" =>  data <= "11111111";  -- 1D48 = FF
      when "1110101001001" =>  data <= "11111111";  -- 1D49 = FF
      when "1110101001010" =>  data <= "11111111";  -- 1D4A = FF
      when "1110101001011" =>  data <= "11111111";  -- 1D4B = FF
      when "1110101001100" =>  data <= "11111111";  -- 1D4C = FF
      when "1110101001101" =>  data <= "11111111";  -- 1D4D = FF
      when "1110101001110" =>  data <= "11111111";  -- 1D4E = FF
      when "1110101001111" =>  data <= "11111111";  -- 1D4F = FF
      when "1110101010000" =>  data <= "11111111";  -- 1D50 = FF
      when "1110101010001" =>  data <= "11111111";  -- 1D51 = FF
      when "1110101010010" =>  data <= "11111111";  -- 1D52 = FF
      when "1110101010011" =>  data <= "11111111";  -- 1D53 = FF
      when "1110101010100" =>  data <= "11111111";  -- 1D54 = FF
      when "1110101010101" =>  data <= "11111111";  -- 1D55 = FF
      when "1110101010110" =>  data <= "11111111";  -- 1D56 = FF
      when "1110101010111" =>  data <= "11111111";  -- 1D57 = FF
      when "1110101011000" =>  data <= "11111111";  -- 1D58 = FF
      when "1110101011001" =>  data <= "11111111";  -- 1D59 = FF
      when "1110101011010" =>  data <= "11111111";  -- 1D5A = FF
      when "1110101011011" =>  data <= "11111111";  -- 1D5B = FF
      when "1110101011100" =>  data <= "11111111";  -- 1D5C = FF
      when "1110101011101" =>  data <= "11111111";  -- 1D5D = FF
      when "1110101011110" =>  data <= "11111111";  -- 1D5E = FF
      when "1110101011111" =>  data <= "11111111";  -- 1D5F = FF
      when "1110101100000" =>  data <= "11111111";  -- 1D60 = FF
      when "1110101100001" =>  data <= "11111111";  -- 1D61 = FF
      when "1110101100010" =>  data <= "11111111";  -- 1D62 = FF
      when "1110101100011" =>  data <= "11111111";  -- 1D63 = FF
      when "1110101100100" =>  data <= "11111111";  -- 1D64 = FF
      when "1110101100101" =>  data <= "11111111";  -- 1D65 = FF
      when "1110101100110" =>  data <= "11111111";  -- 1D66 = FF
      when "1110101100111" =>  data <= "11111111";  -- 1D67 = FF
      when "1110101101000" =>  data <= "11111111";  -- 1D68 = FF
      when "1110101101001" =>  data <= "11111111";  -- 1D69 = FF
      when "1110101101010" =>  data <= "11111111";  -- 1D6A = FF
      when "1110101101011" =>  data <= "11111111";  -- 1D6B = FF
      when "1110101101100" =>  data <= "11111111";  -- 1D6C = FF
      when "1110101101101" =>  data <= "11111111";  -- 1D6D = FF
      when "1110101101110" =>  data <= "11111111";  -- 1D6E = FF
      when "1110101101111" =>  data <= "11111111";  -- 1D6F = FF
      when "1110101110000" =>  data <= "11111111";  -- 1D70 = FF
      when "1110101110001" =>  data <= "11111111";  -- 1D71 = FF
      when "1110101110010" =>  data <= "11111111";  -- 1D72 = FF
      when "1110101110011" =>  data <= "11111111";  -- 1D73 = FF
      when "1110101110100" =>  data <= "11111111";  -- 1D74 = FF
      when "1110101110101" =>  data <= "11111111";  -- 1D75 = FF
      when "1110101110110" =>  data <= "11111111";  -- 1D76 = FF
      when "1110101110111" =>  data <= "11111111";  -- 1D77 = FF
      when "1110101111000" =>  data <= "11111111";  -- 1D78 = FF
      when "1110101111001" =>  data <= "11111111";  -- 1D79 = FF
      when "1110101111010" =>  data <= "11111111";  -- 1D7A = FF
      when "1110101111011" =>  data <= "11111111";  -- 1D7B = FF
      when "1110101111100" =>  data <= "11111111";  -- 1D7C = FF
      when "1110101111101" =>  data <= "11111111";  -- 1D7D = FF
      when "1110101111110" =>  data <= "11111111";  -- 1D7E = FF
      when "1110101111111" =>  data <= "11111111";  -- 1D7F = FF
      when "1110110000000" =>  data <= "11111111";  -- 1D80 = FF
      when "1110110000001" =>  data <= "11111111";  -- 1D81 = FF
      when "1110110000010" =>  data <= "11111111";  -- 1D82 = FF
      when "1110110000011" =>  data <= "11111111";  -- 1D83 = FF
      when "1110110000100" =>  data <= "11111111";  -- 1D84 = FF
      when "1110110000101" =>  data <= "11111111";  -- 1D85 = FF
      when "1110110000110" =>  data <= "11111111";  -- 1D86 = FF
      when "1110110000111" =>  data <= "11111111";  -- 1D87 = FF
      when "1110110001000" =>  data <= "11111111";  -- 1D88 = FF
      when "1110110001001" =>  data <= "11111111";  -- 1D89 = FF
      when "1110110001010" =>  data <= "11111111";  -- 1D8A = FF
      when "1110110001011" =>  data <= "11111111";  -- 1D8B = FF
      when "1110110001100" =>  data <= "11111111";  -- 1D8C = FF
      when "1110110001101" =>  data <= "11111111";  -- 1D8D = FF
      when "1110110001110" =>  data <= "11111111";  -- 1D8E = FF
      when "1110110001111" =>  data <= "11111111";  -- 1D8F = FF
      when "1110110010000" =>  data <= "11111111";  -- 1D90 = FF
      when "1110110010001" =>  data <= "11111111";  -- 1D91 = FF
      when "1110110010010" =>  data <= "11111111";  -- 1D92 = FF
      when "1110110010011" =>  data <= "11111111";  -- 1D93 = FF
      when "1110110010100" =>  data <= "11111111";  -- 1D94 = FF
      when "1110110010101" =>  data <= "11111111";  -- 1D95 = FF
      when "1110110010110" =>  data <= "11111111";  -- 1D96 = FF
      when "1110110010111" =>  data <= "11111111";  -- 1D97 = FF
      when "1110110011000" =>  data <= "11111111";  -- 1D98 = FF
      when "1110110011001" =>  data <= "11111111";  -- 1D99 = FF
      when "1110110011010" =>  data <= "11111111";  -- 1D9A = FF
      when "1110110011011" =>  data <= "11111111";  -- 1D9B = FF
      when "1110110011100" =>  data <= "11111111";  -- 1D9C = FF
      when "1110110011101" =>  data <= "11111111";  -- 1D9D = FF
      when "1110110011110" =>  data <= "11111111";  -- 1D9E = FF
      when "1110110011111" =>  data <= "11111111";  -- 1D9F = FF
      when "1110110100000" =>  data <= "11111111";  -- 1DA0 = FF
      when "1110110100001" =>  data <= "11111111";  -- 1DA1 = FF
      when "1110110100010" =>  data <= "11111111";  -- 1DA2 = FF
      when "1110110100011" =>  data <= "11111111";  -- 1DA3 = FF
      when "1110110100100" =>  data <= "11111111";  -- 1DA4 = FF
      when "1110110100101" =>  data <= "11111111";  -- 1DA5 = FF
      when "1110110100110" =>  data <= "11111111";  -- 1DA6 = FF
      when "1110110100111" =>  data <= "11111111";  -- 1DA7 = FF
      when "1110110101000" =>  data <= "11111111";  -- 1DA8 = FF
      when "1110110101001" =>  data <= "11111111";  -- 1DA9 = FF
      when "1110110101010" =>  data <= "11111111";  -- 1DAA = FF
      when "1110110101011" =>  data <= "11111111";  -- 1DAB = FF
      when "1110110101100" =>  data <= "11111111";  -- 1DAC = FF
      when "1110110101101" =>  data <= "11111111";  -- 1DAD = FF
      when "1110110101110" =>  data <= "11111111";  -- 1DAE = FF
      when "1110110101111" =>  data <= "11111111";  -- 1DAF = FF
      when "1110110110000" =>  data <= "11111111";  -- 1DB0 = FF
      when "1110110110001" =>  data <= "11111111";  -- 1DB1 = FF
      when "1110110110010" =>  data <= "11111111";  -- 1DB2 = FF
      when "1110110110011" =>  data <= "11111111";  -- 1DB3 = FF
      when "1110110110100" =>  data <= "11111111";  -- 1DB4 = FF
      when "1110110110101" =>  data <= "11111111";  -- 1DB5 = FF
      when "1110110110110" =>  data <= "11111111";  -- 1DB6 = FF
      when "1110110110111" =>  data <= "11111111";  -- 1DB7 = FF
      when "1110110111000" =>  data <= "11111111";  -- 1DB8 = FF
      when "1110110111001" =>  data <= "11111111";  -- 1DB9 = FF
      when "1110110111010" =>  data <= "11111111";  -- 1DBA = FF
      when "1110110111011" =>  data <= "11111111";  -- 1DBB = FF
      when "1110110111100" =>  data <= "11111111";  -- 1DBC = FF
      when "1110110111101" =>  data <= "11111111";  -- 1DBD = FF
      when "1110110111110" =>  data <= "11111111";  -- 1DBE = FF
      when "1110110111111" =>  data <= "11111111";  -- 1DBF = FF
      when "1110111000000" =>  data <= "11111111";  -- 1DC0 = FF
      when "1110111000001" =>  data <= "11111111";  -- 1DC1 = FF
      when "1110111000010" =>  data <= "11111111";  -- 1DC2 = FF
      when "1110111000011" =>  data <= "11111111";  -- 1DC3 = FF
      when "1110111000100" =>  data <= "11111111";  -- 1DC4 = FF
      when "1110111000101" =>  data <= "11111111";  -- 1DC5 = FF
      when "1110111000110" =>  data <= "11111111";  -- 1DC6 = FF
      when "1110111000111" =>  data <= "11111111";  -- 1DC7 = FF
      when "1110111001000" =>  data <= "11111111";  -- 1DC8 = FF
      when "1110111001001" =>  data <= "11111111";  -- 1DC9 = FF
      when "1110111001010" =>  data <= "11111111";  -- 1DCA = FF
      when "1110111001011" =>  data <= "11111111";  -- 1DCB = FF
      when "1110111001100" =>  data <= "11111111";  -- 1DCC = FF
      when "1110111001101" =>  data <= "11111111";  -- 1DCD = FF
      when "1110111001110" =>  data <= "11111111";  -- 1DCE = FF
      when "1110111001111" =>  data <= "11111111";  -- 1DCF = FF
      when "1110111010000" =>  data <= "11111111";  -- 1DD0 = FF
      when "1110111010001" =>  data <= "11111111";  -- 1DD1 = FF
      when "1110111010010" =>  data <= "11111111";  -- 1DD2 = FF
      when "1110111010011" =>  data <= "11111111";  -- 1DD3 = FF
      when "1110111010100" =>  data <= "11111111";  -- 1DD4 = FF
      when "1110111010101" =>  data <= "11111111";  -- 1DD5 = FF
      when "1110111010110" =>  data <= "11111111";  -- 1DD6 = FF
      when "1110111010111" =>  data <= "11111111";  -- 1DD7 = FF
      when "1110111011000" =>  data <= "11111111";  -- 1DD8 = FF
      when "1110111011001" =>  data <= "11111111";  -- 1DD9 = FF
      when "1110111011010" =>  data <= "11111111";  -- 1DDA = FF
      when "1110111011011" =>  data <= "11111111";  -- 1DDB = FF
      when "1110111011100" =>  data <= "11111111";  -- 1DDC = FF
      when "1110111011101" =>  data <= "11111111";  -- 1DDD = FF
      when "1110111011110" =>  data <= "11111111";  -- 1DDE = FF
      when "1110111011111" =>  data <= "11111111";  -- 1DDF = FF
      when "1110111100000" =>  data <= "11111111";  -- 1DE0 = FF
      when "1110111100001" =>  data <= "11111111";  -- 1DE1 = FF
      when "1110111100010" =>  data <= "11111111";  -- 1DE2 = FF
      when "1110111100011" =>  data <= "11111111";  -- 1DE3 = FF
      when "1110111100100" =>  data <= "11111111";  -- 1DE4 = FF
      when "1110111100101" =>  data <= "11111111";  -- 1DE5 = FF
      when "1110111100110" =>  data <= "11111111";  -- 1DE6 = FF
      when "1110111100111" =>  data <= "11111111";  -- 1DE7 = FF
      when "1110111101000" =>  data <= "11111111";  -- 1DE8 = FF
      when "1110111101001" =>  data <= "11111111";  -- 1DE9 = FF
      when "1110111101010" =>  data <= "11111111";  -- 1DEA = FF
      when "1110111101011" =>  data <= "11111111";  -- 1DEB = FF
      when "1110111101100" =>  data <= "11111111";  -- 1DEC = FF
      when "1110111101101" =>  data <= "11111111";  -- 1DED = FF
      when "1110111101110" =>  data <= "11111111";  -- 1DEE = FF
      when "1110111101111" =>  data <= "11111111";  -- 1DEF = FF
      when "1110111110000" =>  data <= "11111111";  -- 1DF0 = FF
      when "1110111110001" =>  data <= "11111111";  -- 1DF1 = FF
      when "1110111110010" =>  data <= "11111111";  -- 1DF2 = FF
      when "1110111110011" =>  data <= "11111111";  -- 1DF3 = FF
      when "1110111110100" =>  data <= "11111111";  -- 1DF4 = FF
      when "1110111110101" =>  data <= "11111111";  -- 1DF5 = FF
      when "1110111110110" =>  data <= "11111111";  -- 1DF6 = FF
      when "1110111110111" =>  data <= "11111111";  -- 1DF7 = FF
      when "1110111111000" =>  data <= "11111111";  -- 1DF8 = FF
      when "1110111111001" =>  data <= "11111111";  -- 1DF9 = FF
      when "1110111111010" =>  data <= "11111111";  -- 1DFA = FF
      when "1110111111011" =>  data <= "11111111";  -- 1DFB = FF
      when "1110111111100" =>  data <= "11111111";  -- 1DFC = FF
      when "1110111111101" =>  data <= "11111111";  -- 1DFD = FF
      when "1110111111110" =>  data <= "11111111";  -- 1DFE = FF
      when "1110111111111" =>  data <= "11111111";  -- 1DFF = FF
      when "1111000000000" =>  data <= "11111111";  -- 1E00 = FF
      when "1111000000001" =>  data <= "11111111";  -- 1E01 = FF
      when "1111000000010" =>  data <= "11111111";  -- 1E02 = FF
      when "1111000000011" =>  data <= "11111111";  -- 1E03 = FF
      when "1111000000100" =>  data <= "11111111";  -- 1E04 = FF
      when "1111000000101" =>  data <= "11111111";  -- 1E05 = FF
      when "1111000000110" =>  data <= "11111111";  -- 1E06 = FF
      when "1111000000111" =>  data <= "11111111";  -- 1E07 = FF
      when "1111000001000" =>  data <= "11111111";  -- 1E08 = FF
      when "1111000001001" =>  data <= "11111111";  -- 1E09 = FF
      when "1111000001010" =>  data <= "11111111";  -- 1E0A = FF
      when "1111000001011" =>  data <= "11111111";  -- 1E0B = FF
      when "1111000001100" =>  data <= "11111111";  -- 1E0C = FF
      when "1111000001101" =>  data <= "11111111";  -- 1E0D = FF
      when "1111000001110" =>  data <= "11111111";  -- 1E0E = FF
      when "1111000001111" =>  data <= "11111111";  -- 1E0F = FF
      when "1111000010000" =>  data <= "11111111";  -- 1E10 = FF
      when "1111000010001" =>  data <= "11111111";  -- 1E11 = FF
      when "1111000010010" =>  data <= "11111111";  -- 1E12 = FF
      when "1111000010011" =>  data <= "11111111";  -- 1E13 = FF
      when "1111000010100" =>  data <= "11111111";  -- 1E14 = FF
      when "1111000010101" =>  data <= "11111111";  -- 1E15 = FF
      when "1111000010110" =>  data <= "11111111";  -- 1E16 = FF
      when "1111000010111" =>  data <= "11111111";  -- 1E17 = FF
      when "1111000011000" =>  data <= "11111111";  -- 1E18 = FF
      when "1111000011001" =>  data <= "11111111";  -- 1E19 = FF
      when "1111000011010" =>  data <= "11111111";  -- 1E1A = FF
      when "1111000011011" =>  data <= "11111111";  -- 1E1B = FF
      when "1111000011100" =>  data <= "11111111";  -- 1E1C = FF
      when "1111000011101" =>  data <= "11111111";  -- 1E1D = FF
      when "1111000011110" =>  data <= "11111111";  -- 1E1E = FF
      when "1111000011111" =>  data <= "11111111";  -- 1E1F = FF
      when "1111000100000" =>  data <= "11111111";  -- 1E20 = FF
      when "1111000100001" =>  data <= "11111111";  -- 1E21 = FF
      when "1111000100010" =>  data <= "11111111";  -- 1E22 = FF
      when "1111000100011" =>  data <= "11111111";  -- 1E23 = FF
      when "1111000100100" =>  data <= "11111111";  -- 1E24 = FF
      when "1111000100101" =>  data <= "11111111";  -- 1E25 = FF
      when "1111000100110" =>  data <= "11111111";  -- 1E26 = FF
      when "1111000100111" =>  data <= "11111111";  -- 1E27 = FF
      when "1111000101000" =>  data <= "11111111";  -- 1E28 = FF
      when "1111000101001" =>  data <= "11111111";  -- 1E29 = FF
      when "1111000101010" =>  data <= "11111111";  -- 1E2A = FF
      when "1111000101011" =>  data <= "11111111";  -- 1E2B = FF
      when "1111000101100" =>  data <= "11111111";  -- 1E2C = FF
      when "1111000101101" =>  data <= "11111111";  -- 1E2D = FF
      when "1111000101110" =>  data <= "11111111";  -- 1E2E = FF
      when "1111000101111" =>  data <= "11111111";  -- 1E2F = FF
      when "1111000110000" =>  data <= "11111111";  -- 1E30 = FF
      when "1111000110001" =>  data <= "11111111";  -- 1E31 = FF
      when "1111000110010" =>  data <= "11111111";  -- 1E32 = FF
      when "1111000110011" =>  data <= "11111111";  -- 1E33 = FF
      when "1111000110100" =>  data <= "11111111";  -- 1E34 = FF
      when "1111000110101" =>  data <= "11111111";  -- 1E35 = FF
      when "1111000110110" =>  data <= "11111111";  -- 1E36 = FF
      when "1111000110111" =>  data <= "11111111";  -- 1E37 = FF
      when "1111000111000" =>  data <= "11111111";  -- 1E38 = FF
      when "1111000111001" =>  data <= "11111111";  -- 1E39 = FF
      when "1111000111010" =>  data <= "11111111";  -- 1E3A = FF
      when "1111000111011" =>  data <= "11111111";  -- 1E3B = FF
      when "1111000111100" =>  data <= "11111111";  -- 1E3C = FF
      when "1111000111101" =>  data <= "11111111";  -- 1E3D = FF
      when "1111000111110" =>  data <= "11111111";  -- 1E3E = FF
      when "1111000111111" =>  data <= "11111111";  -- 1E3F = FF
      when "1111001000000" =>  data <= "11111111";  -- 1E40 = FF
      when "1111001000001" =>  data <= "11111111";  -- 1E41 = FF
      when "1111001000010" =>  data <= "11111111";  -- 1E42 = FF
      when "1111001000011" =>  data <= "11111111";  -- 1E43 = FF
      when "1111001000100" =>  data <= "11111111";  -- 1E44 = FF
      when "1111001000101" =>  data <= "11111111";  -- 1E45 = FF
      when "1111001000110" =>  data <= "11111111";  -- 1E46 = FF
      when "1111001000111" =>  data <= "11111111";  -- 1E47 = FF
      when "1111001001000" =>  data <= "11111111";  -- 1E48 = FF
      when "1111001001001" =>  data <= "11111111";  -- 1E49 = FF
      when "1111001001010" =>  data <= "11111111";  -- 1E4A = FF
      when "1111001001011" =>  data <= "11111111";  -- 1E4B = FF
      when "1111001001100" =>  data <= "11111111";  -- 1E4C = FF
      when "1111001001101" =>  data <= "11111111";  -- 1E4D = FF
      when "1111001001110" =>  data <= "11111111";  -- 1E4E = FF
      when "1111001001111" =>  data <= "11111111";  -- 1E4F = FF
      when "1111001010000" =>  data <= "11111111";  -- 1E50 = FF
      when "1111001010001" =>  data <= "11111111";  -- 1E51 = FF
      when "1111001010010" =>  data <= "11111111";  -- 1E52 = FF
      when "1111001010011" =>  data <= "11111111";  -- 1E53 = FF
      when "1111001010100" =>  data <= "11111111";  -- 1E54 = FF
      when "1111001010101" =>  data <= "11111111";  -- 1E55 = FF
      when "1111001010110" =>  data <= "11111111";  -- 1E56 = FF
      when "1111001010111" =>  data <= "11111111";  -- 1E57 = FF
      when "1111001011000" =>  data <= "11111111";  -- 1E58 = FF
      when "1111001011001" =>  data <= "11111111";  -- 1E59 = FF
      when "1111001011010" =>  data <= "11111111";  -- 1E5A = FF
      when "1111001011011" =>  data <= "11111111";  -- 1E5B = FF
      when "1111001011100" =>  data <= "11111111";  -- 1E5C = FF
      when "1111001011101" =>  data <= "11111111";  -- 1E5D = FF
      when "1111001011110" =>  data <= "11111111";  -- 1E5E = FF
      when "1111001011111" =>  data <= "11111111";  -- 1E5F = FF
      when "1111001100000" =>  data <= "11111111";  -- 1E60 = FF
      when "1111001100001" =>  data <= "11111111";  -- 1E61 = FF
      when "1111001100010" =>  data <= "11111111";  -- 1E62 = FF
      when "1111001100011" =>  data <= "11111111";  -- 1E63 = FF
      when "1111001100100" =>  data <= "11111111";  -- 1E64 = FF
      when "1111001100101" =>  data <= "11111111";  -- 1E65 = FF
      when "1111001100110" =>  data <= "11111111";  -- 1E66 = FF
      when "1111001100111" =>  data <= "11111111";  -- 1E67 = FF
      when "1111001101000" =>  data <= "11111111";  -- 1E68 = FF
      when "1111001101001" =>  data <= "11111111";  -- 1E69 = FF
      when "1111001101010" =>  data <= "11111111";  -- 1E6A = FF
      when "1111001101011" =>  data <= "11111111";  -- 1E6B = FF
      when "1111001101100" =>  data <= "11111111";  -- 1E6C = FF
      when "1111001101101" =>  data <= "11111111";  -- 1E6D = FF
      when "1111001101110" =>  data <= "11111111";  -- 1E6E = FF
      when "1111001101111" =>  data <= "11111111";  -- 1E6F = FF
      when "1111001110000" =>  data <= "11111111";  -- 1E70 = FF
      when "1111001110001" =>  data <= "11111111";  -- 1E71 = FF
      when "1111001110010" =>  data <= "11111111";  -- 1E72 = FF
      when "1111001110011" =>  data <= "11111111";  -- 1E73 = FF
      when "1111001110100" =>  data <= "11111111";  -- 1E74 = FF
      when "1111001110101" =>  data <= "11111111";  -- 1E75 = FF
      when "1111001110110" =>  data <= "11111111";  -- 1E76 = FF
      when "1111001110111" =>  data <= "11111111";  -- 1E77 = FF
      when "1111001111000" =>  data <= "11111111";  -- 1E78 = FF
      when "1111001111001" =>  data <= "11111111";  -- 1E79 = FF
      when "1111001111010" =>  data <= "11111111";  -- 1E7A = FF
      when "1111001111011" =>  data <= "11111111";  -- 1E7B = FF
      when "1111001111100" =>  data <= "11111111";  -- 1E7C = FF
      when "1111001111101" =>  data <= "11111111";  -- 1E7D = FF
      when "1111001111110" =>  data <= "11111111";  -- 1E7E = FF
      when "1111001111111" =>  data <= "11111111";  -- 1E7F = FF
      when "1111010000000" =>  data <= "11111111";  -- 1E80 = FF
      when "1111010000001" =>  data <= "11111111";  -- 1E81 = FF
      when "1111010000010" =>  data <= "11111111";  -- 1E82 = FF
      when "1111010000011" =>  data <= "11111111";  -- 1E83 = FF
      when "1111010000100" =>  data <= "11111111";  -- 1E84 = FF
      when "1111010000101" =>  data <= "11111111";  -- 1E85 = FF
      when "1111010000110" =>  data <= "11111111";  -- 1E86 = FF
      when "1111010000111" =>  data <= "11111111";  -- 1E87 = FF
      when "1111010001000" =>  data <= "11111111";  -- 1E88 = FF
      when "1111010001001" =>  data <= "11111111";  -- 1E89 = FF
      when "1111010001010" =>  data <= "11111111";  -- 1E8A = FF
      when "1111010001011" =>  data <= "11111111";  -- 1E8B = FF
      when "1111010001100" =>  data <= "11111111";  -- 1E8C = FF
      when "1111010001101" =>  data <= "11111111";  -- 1E8D = FF
      when "1111010001110" =>  data <= "11111111";  -- 1E8E = FF
      when "1111010001111" =>  data <= "11111111";  -- 1E8F = FF
      when "1111010010000" =>  data <= "11111111";  -- 1E90 = FF
      when "1111010010001" =>  data <= "11111111";  -- 1E91 = FF
      when "1111010010010" =>  data <= "11111111";  -- 1E92 = FF
      when "1111010010011" =>  data <= "11111111";  -- 1E93 = FF
      when "1111010010100" =>  data <= "11111111";  -- 1E94 = FF
      when "1111010010101" =>  data <= "11111111";  -- 1E95 = FF
      when "1111010010110" =>  data <= "11111111";  -- 1E96 = FF
      when "1111010010111" =>  data <= "11111111";  -- 1E97 = FF
      when "1111010011000" =>  data <= "11111111";  -- 1E98 = FF
      when "1111010011001" =>  data <= "11111111";  -- 1E99 = FF
      when "1111010011010" =>  data <= "11111111";  -- 1E9A = FF
      when "1111010011011" =>  data <= "11111111";  -- 1E9B = FF
      when "1111010011100" =>  data <= "11111111";  -- 1E9C = FF
      when "1111010011101" =>  data <= "11111111";  -- 1E9D = FF
      when "1111010011110" =>  data <= "11111111";  -- 1E9E = FF
      when "1111010011111" =>  data <= "11111111";  -- 1E9F = FF
      when "1111010100000" =>  data <= "11111111";  -- 1EA0 = FF
      when "1111010100001" =>  data <= "11111111";  -- 1EA1 = FF
      when "1111010100010" =>  data <= "11111111";  -- 1EA2 = FF
      when "1111010100011" =>  data <= "11111111";  -- 1EA3 = FF
      when "1111010100100" =>  data <= "11111111";  -- 1EA4 = FF
      when "1111010100101" =>  data <= "11111111";  -- 1EA5 = FF
      when "1111010100110" =>  data <= "11111111";  -- 1EA6 = FF
      when "1111010100111" =>  data <= "11111111";  -- 1EA7 = FF
      when "1111010101000" =>  data <= "11111111";  -- 1EA8 = FF
      when "1111010101001" =>  data <= "11111111";  -- 1EA9 = FF
      when "1111010101010" =>  data <= "11111111";  -- 1EAA = FF
      when "1111010101011" =>  data <= "11111111";  -- 1EAB = FF
      when "1111010101100" =>  data <= "11111111";  -- 1EAC = FF
      when "1111010101101" =>  data <= "11111111";  -- 1EAD = FF
      when "1111010101110" =>  data <= "11111111";  -- 1EAE = FF
      when "1111010101111" =>  data <= "11111111";  -- 1EAF = FF
      when "1111010110000" =>  data <= "11111111";  -- 1EB0 = FF
      when "1111010110001" =>  data <= "11111111";  -- 1EB1 = FF
      when "1111010110010" =>  data <= "11111111";  -- 1EB2 = FF
      when "1111010110011" =>  data <= "11111111";  -- 1EB3 = FF
      when "1111010110100" =>  data <= "11111111";  -- 1EB4 = FF
      when "1111010110101" =>  data <= "11111111";  -- 1EB5 = FF
      when "1111010110110" =>  data <= "11111111";  -- 1EB6 = FF
      when "1111010110111" =>  data <= "11111111";  -- 1EB7 = FF
      when "1111010111000" =>  data <= "11111111";  -- 1EB8 = FF
      when "1111010111001" =>  data <= "11111111";  -- 1EB9 = FF
      when "1111010111010" =>  data <= "11111111";  -- 1EBA = FF
      when "1111010111011" =>  data <= "11111111";  -- 1EBB = FF
      when "1111010111100" =>  data <= "11111111";  -- 1EBC = FF
      when "1111010111101" =>  data <= "11111111";  -- 1EBD = FF
      when "1111010111110" =>  data <= "11111111";  -- 1EBE = FF
      when "1111010111111" =>  data <= "11111111";  -- 1EBF = FF
      when "1111011000000" =>  data <= "11111111";  -- 1EC0 = FF
      when "1111011000001" =>  data <= "11111111";  -- 1EC1 = FF
      when "1111011000010" =>  data <= "11111111";  -- 1EC2 = FF
      when "1111011000011" =>  data <= "11111111";  -- 1EC3 = FF
      when "1111011000100" =>  data <= "11111111";  -- 1EC4 = FF
      when "1111011000101" =>  data <= "11111111";  -- 1EC5 = FF
      when "1111011000110" =>  data <= "11111111";  -- 1EC6 = FF
      when "1111011000111" =>  data <= "11111111";  -- 1EC7 = FF
      when "1111011001000" =>  data <= "11111111";  -- 1EC8 = FF
      when "1111011001001" =>  data <= "11111111";  -- 1EC9 = FF
      when "1111011001010" =>  data <= "11111111";  -- 1ECA = FF
      when "1111011001011" =>  data <= "11111111";  -- 1ECB = FF
      when "1111011001100" =>  data <= "11111111";  -- 1ECC = FF
      when "1111011001101" =>  data <= "11111111";  -- 1ECD = FF
      when "1111011001110" =>  data <= "11111111";  -- 1ECE = FF
      when "1111011001111" =>  data <= "11111111";  -- 1ECF = FF
      when "1111011010000" =>  data <= "11111111";  -- 1ED0 = FF
      when "1111011010001" =>  data <= "11111111";  -- 1ED1 = FF
      when "1111011010010" =>  data <= "11111111";  -- 1ED2 = FF
      when "1111011010011" =>  data <= "11111111";  -- 1ED3 = FF
      when "1111011010100" =>  data <= "11111111";  -- 1ED4 = FF
      when "1111011010101" =>  data <= "11111111";  -- 1ED5 = FF
      when "1111011010110" =>  data <= "11111111";  -- 1ED6 = FF
      when "1111011010111" =>  data <= "11111111";  -- 1ED7 = FF
      when "1111011011000" =>  data <= "11111111";  -- 1ED8 = FF
      when "1111011011001" =>  data <= "11111111";  -- 1ED9 = FF
      when "1111011011010" =>  data <= "11111111";  -- 1EDA = FF
      when "1111011011011" =>  data <= "11111111";  -- 1EDB = FF
      when "1111011011100" =>  data <= "11111111";  -- 1EDC = FF
      when "1111011011101" =>  data <= "11111111";  -- 1EDD = FF
      when "1111011011110" =>  data <= "11111111";  -- 1EDE = FF
      when "1111011011111" =>  data <= "11111111";  -- 1EDF = FF
      when "1111011100000" =>  data <= "11111111";  -- 1EE0 = FF
      when "1111011100001" =>  data <= "11111111";  -- 1EE1 = FF
      when "1111011100010" =>  data <= "11111111";  -- 1EE2 = FF
      when "1111011100011" =>  data <= "11111111";  -- 1EE3 = FF
      when "1111011100100" =>  data <= "11111111";  -- 1EE4 = FF
      when "1111011100101" =>  data <= "11111111";  -- 1EE5 = FF
      when "1111011100110" =>  data <= "11111111";  -- 1EE6 = FF
      when "1111011100111" =>  data <= "11111111";  -- 1EE7 = FF
      when "1111011101000" =>  data <= "11111111";  -- 1EE8 = FF
      when "1111011101001" =>  data <= "11111111";  -- 1EE9 = FF
      when "1111011101010" =>  data <= "11111111";  -- 1EEA = FF
      when "1111011101011" =>  data <= "11111111";  -- 1EEB = FF
      when "1111011101100" =>  data <= "11111111";  -- 1EEC = FF
      when "1111011101101" =>  data <= "11111111";  -- 1EED = FF
      when "1111011101110" =>  data <= "11111111";  -- 1EEE = FF
      when "1111011101111" =>  data <= "11111111";  -- 1EEF = FF
      when "1111011110000" =>  data <= "11111111";  -- 1EF0 = FF
      when "1111011110001" =>  data <= "11111111";  -- 1EF1 = FF
      when "1111011110010" =>  data <= "11111111";  -- 1EF2 = FF
      when "1111011110011" =>  data <= "11111111";  -- 1EF3 = FF
      when "1111011110100" =>  data <= "11111111";  -- 1EF4 = FF
      when "1111011110101" =>  data <= "11111111";  -- 1EF5 = FF
      when "1111011110110" =>  data <= "11111111";  -- 1EF6 = FF
      when "1111011110111" =>  data <= "11111111";  -- 1EF7 = FF
      when "1111011111000" =>  data <= "11111111";  -- 1EF8 = FF
      when "1111011111001" =>  data <= "11111111";  -- 1EF9 = FF
      when "1111011111010" =>  data <= "11111111";  -- 1EFA = FF
      when "1111011111011" =>  data <= "11111111";  -- 1EFB = FF
      when "1111011111100" =>  data <= "11111111";  -- 1EFC = FF
      when "1111011111101" =>  data <= "11111111";  -- 1EFD = FF
      when "1111011111110" =>  data <= "11111111";  -- 1EFE = FF
      when "1111011111111" =>  data <= "11111111";  -- 1EFF = FF
      when "1111100000000" =>  data <= "11111111";  -- 1F00 = FF
      when "1111100000001" =>  data <= "11111111";  -- 1F01 = FF
      when "1111100000010" =>  data <= "11111111";  -- 1F02 = FF
      when "1111100000011" =>  data <= "11111111";  -- 1F03 = FF
      when "1111100000100" =>  data <= "11111111";  -- 1F04 = FF
      when "1111100000101" =>  data <= "11111111";  -- 1F05 = FF
      when "1111100000110" =>  data <= "11111111";  -- 1F06 = FF
      when "1111100000111" =>  data <= "11111111";  -- 1F07 = FF
      when "1111100001000" =>  data <= "11111111";  -- 1F08 = FF
      when "1111100001001" =>  data <= "11111111";  -- 1F09 = FF
      when "1111100001010" =>  data <= "11111111";  -- 1F0A = FF
      when "1111100001011" =>  data <= "11111111";  -- 1F0B = FF
      when "1111100001100" =>  data <= "11111111";  -- 1F0C = FF
      when "1111100001101" =>  data <= "11111111";  -- 1F0D = FF
      when "1111100001110" =>  data <= "11111111";  -- 1F0E = FF
      when "1111100001111" =>  data <= "11111111";  -- 1F0F = FF
      when "1111100010000" =>  data <= "11111111";  -- 1F10 = FF
      when "1111100010001" =>  data <= "11111111";  -- 1F11 = FF
      when "1111100010010" =>  data <= "11111111";  -- 1F12 = FF
      when "1111100010011" =>  data <= "11111111";  -- 1F13 = FF
      when "1111100010100" =>  data <= "11111111";  -- 1F14 = FF
      when "1111100010101" =>  data <= "11111111";  -- 1F15 = FF
      when "1111100010110" =>  data <= "11111111";  -- 1F16 = FF
      when "1111100010111" =>  data <= "11111111";  -- 1F17 = FF
      when "1111100011000" =>  data <= "11111111";  -- 1F18 = FF
      when "1111100011001" =>  data <= "11111111";  -- 1F19 = FF
      when "1111100011010" =>  data <= "11111111";  -- 1F1A = FF
      when "1111100011011" =>  data <= "11111111";  -- 1F1B = FF
      when "1111100011100" =>  data <= "11111111";  -- 1F1C = FF
      when "1111100011101" =>  data <= "11111111";  -- 1F1D = FF
      when "1111100011110" =>  data <= "11111111";  -- 1F1E = FF
      when "1111100011111" =>  data <= "11111111";  -- 1F1F = FF
      when "1111100100000" =>  data <= "11111111";  -- 1F20 = FF
      when "1111100100001" =>  data <= "11111111";  -- 1F21 = FF
      when "1111100100010" =>  data <= "11111111";  -- 1F22 = FF
      when "1111100100011" =>  data <= "11111111";  -- 1F23 = FF
      when "1111100100100" =>  data <= "11111111";  -- 1F24 = FF
      when "1111100100101" =>  data <= "11111111";  -- 1F25 = FF
      when "1111100100110" =>  data <= "11111111";  -- 1F26 = FF
      when "1111100100111" =>  data <= "11111111";  -- 1F27 = FF
      when "1111100101000" =>  data <= "11111111";  -- 1F28 = FF
      when "1111100101001" =>  data <= "11111111";  -- 1F29 = FF
      when "1111100101010" =>  data <= "11111111";  -- 1F2A = FF
      when "1111100101011" =>  data <= "11111111";  -- 1F2B = FF
      when "1111100101100" =>  data <= "11111111";  -- 1F2C = FF
      when "1111100101101" =>  data <= "11111111";  -- 1F2D = FF
      when "1111100101110" =>  data <= "11111111";  -- 1F2E = FF
      when "1111100101111" =>  data <= "11111111";  -- 1F2F = FF
      when "1111100110000" =>  data <= "11111111";  -- 1F30 = FF
      when "1111100110001" =>  data <= "11111111";  -- 1F31 = FF
      when "1111100110010" =>  data <= "11111111";  -- 1F32 = FF
      when "1111100110011" =>  data <= "11111111";  -- 1F33 = FF
      when "1111100110100" =>  data <= "11111111";  -- 1F34 = FF
      when "1111100110101" =>  data <= "11111111";  -- 1F35 = FF
      when "1111100110110" =>  data <= "11111111";  -- 1F36 = FF
      when "1111100110111" =>  data <= "11111111";  -- 1F37 = FF
      when "1111100111000" =>  data <= "11111111";  -- 1F38 = FF
      when "1111100111001" =>  data <= "11111111";  -- 1F39 = FF
      when "1111100111010" =>  data <= "11111111";  -- 1F3A = FF
      when "1111100111011" =>  data <= "11111111";  -- 1F3B = FF
      when "1111100111100" =>  data <= "11111111";  -- 1F3C = FF
      when "1111100111101" =>  data <= "11111111";  -- 1F3D = FF
      when "1111100111110" =>  data <= "11111111";  -- 1F3E = FF
      when "1111100111111" =>  data <= "11111111";  -- 1F3F = FF
      when "1111101000000" =>  data <= "11111111";  -- 1F40 = FF
      when "1111101000001" =>  data <= "11111111";  -- 1F41 = FF
      when "1111101000010" =>  data <= "11111111";  -- 1F42 = FF
      when "1111101000011" =>  data <= "11111111";  -- 1F43 = FF
      when "1111101000100" =>  data <= "11111111";  -- 1F44 = FF
      when "1111101000101" =>  data <= "11111111";  -- 1F45 = FF
      when "1111101000110" =>  data <= "11111111";  -- 1F46 = FF
      when "1111101000111" =>  data <= "11111111";  -- 1F47 = FF
      when "1111101001000" =>  data <= "11111111";  -- 1F48 = FF
      when "1111101001001" =>  data <= "11111111";  -- 1F49 = FF
      when "1111101001010" =>  data <= "11111111";  -- 1F4A = FF
      when "1111101001011" =>  data <= "11111111";  -- 1F4B = FF
      when "1111101001100" =>  data <= "11111111";  -- 1F4C = FF
      when "1111101001101" =>  data <= "11111111";  -- 1F4D = FF
      when "1111101001110" =>  data <= "11111111";  -- 1F4E = FF
      when "1111101001111" =>  data <= "11111111";  -- 1F4F = FF
      when "1111101010000" =>  data <= "11111111";  -- 1F50 = FF
      when "1111101010001" =>  data <= "11111111";  -- 1F51 = FF
      when "1111101010010" =>  data <= "11111111";  -- 1F52 = FF
      when "1111101010011" =>  data <= "11111111";  -- 1F53 = FF
      when "1111101010100" =>  data <= "11111111";  -- 1F54 = FF
      when "1111101010101" =>  data <= "11111111";  -- 1F55 = FF
      when "1111101010110" =>  data <= "11111111";  -- 1F56 = FF
      when "1111101010111" =>  data <= "11111111";  -- 1F57 = FF
      when "1111101011000" =>  data <= "11111111";  -- 1F58 = FF
      when "1111101011001" =>  data <= "11111111";  -- 1F59 = FF
      when "1111101011010" =>  data <= "11111111";  -- 1F5A = FF
      when "1111101011011" =>  data <= "11111111";  -- 1F5B = FF
      when "1111101011100" =>  data <= "11111111";  -- 1F5C = FF
      when "1111101011101" =>  data <= "11111111";  -- 1F5D = FF
      when "1111101011110" =>  data <= "11111111";  -- 1F5E = FF
      when "1111101011111" =>  data <= "11111111";  -- 1F5F = FF
      when "1111101100000" =>  data <= "11111111";  -- 1F60 = FF
      when "1111101100001" =>  data <= "11111111";  -- 1F61 = FF
      when "1111101100010" =>  data <= "11111111";  -- 1F62 = FF
      when "1111101100011" =>  data <= "11111111";  -- 1F63 = FF
      when "1111101100100" =>  data <= "11111111";  -- 1F64 = FF
      when "1111101100101" =>  data <= "11111111";  -- 1F65 = FF
      when "1111101100110" =>  data <= "11111111";  -- 1F66 = FF
      when "1111101100111" =>  data <= "11111111";  -- 1F67 = FF
      when "1111101101000" =>  data <= "11111111";  -- 1F68 = FF
      when "1111101101001" =>  data <= "11111111";  -- 1F69 = FF
      when "1111101101010" =>  data <= "11111111";  -- 1F6A = FF
      when "1111101101011" =>  data <= "11111111";  -- 1F6B = FF
      when "1111101101100" =>  data <= "11111111";  -- 1F6C = FF
      when "1111101101101" =>  data <= "11111111";  -- 1F6D = FF
      when "1111101101110" =>  data <= "11111111";  -- 1F6E = FF
      when "1111101101111" =>  data <= "11111111";  -- 1F6F = FF
      when "1111101110000" =>  data <= "11111111";  -- 1F70 = FF
      when "1111101110001" =>  data <= "11111111";  -- 1F71 = FF
      when "1111101110010" =>  data <= "11111111";  -- 1F72 = FF
      when "1111101110011" =>  data <= "11111111";  -- 1F73 = FF
      when "1111101110100" =>  data <= "11111111";  -- 1F74 = FF
      when "1111101110101" =>  data <= "11111111";  -- 1F75 = FF
      when "1111101110110" =>  data <= "11111111";  -- 1F76 = FF
      when "1111101110111" =>  data <= "11111111";  -- 1F77 = FF
      when "1111101111000" =>  data <= "11111111";  -- 1F78 = FF
      when "1111101111001" =>  data <= "11111111";  -- 1F79 = FF
      when "1111101111010" =>  data <= "11111111";  -- 1F7A = FF
      when "1111101111011" =>  data <= "11111111";  -- 1F7B = FF
      when "1111101111100" =>  data <= "11111111";  -- 1F7C = FF
      when "1111101111101" =>  data <= "11111111";  -- 1F7D = FF
      when "1111101111110" =>  data <= "11111111";  -- 1F7E = FF
      when "1111101111111" =>  data <= "11111111";  -- 1F7F = FF
      when "1111110000000" =>  data <= "11111111";  -- 1F80 = FF
      when "1111110000001" =>  data <= "11111111";  -- 1F81 = FF
      when "1111110000010" =>  data <= "11111111";  -- 1F82 = FF
      when "1111110000011" =>  data <= "11111111";  -- 1F83 = FF
      when "1111110000100" =>  data <= "11111111";  -- 1F84 = FF
      when "1111110000101" =>  data <= "11111111";  -- 1F85 = FF
      when "1111110000110" =>  data <= "11111111";  -- 1F86 = FF
      when "1111110000111" =>  data <= "11111111";  -- 1F87 = FF
      when "1111110001000" =>  data <= "11111111";  -- 1F88 = FF
      when "1111110001001" =>  data <= "11111111";  -- 1F89 = FF
      when "1111110001010" =>  data <= "11111111";  -- 1F8A = FF
      when "1111110001011" =>  data <= "11111111";  -- 1F8B = FF
      when "1111110001100" =>  data <= "11111111";  -- 1F8C = FF
      when "1111110001101" =>  data <= "11111111";  -- 1F8D = FF
      when "1111110001110" =>  data <= "11111111";  -- 1F8E = FF
      when "1111110001111" =>  data <= "11111111";  -- 1F8F = FF
      when "1111110010000" =>  data <= "11111111";  -- 1F90 = FF
      when "1111110010001" =>  data <= "11111111";  -- 1F91 = FF
      when "1111110010010" =>  data <= "11111111";  -- 1F92 = FF
      when "1111110010011" =>  data <= "11111111";  -- 1F93 = FF
      when "1111110010100" =>  data <= "11111111";  -- 1F94 = FF
      when "1111110010101" =>  data <= "11111111";  -- 1F95 = FF
      when "1111110010110" =>  data <= "11111111";  -- 1F96 = FF
      when "1111110010111" =>  data <= "11111111";  -- 1F97 = FF
      when "1111110011000" =>  data <= "11111111";  -- 1F98 = FF
      when "1111110011001" =>  data <= "11111111";  -- 1F99 = FF
      when "1111110011010" =>  data <= "11111111";  -- 1F9A = FF
      when "1111110011011" =>  data <= "11111111";  -- 1F9B = FF
      when "1111110011100" =>  data <= "11111111";  -- 1F9C = FF
      when "1111110011101" =>  data <= "11111111";  -- 1F9D = FF
      when "1111110011110" =>  data <= "11111111";  -- 1F9E = FF
      when "1111110011111" =>  data <= "11111111";  -- 1F9F = FF
      when "1111110100000" =>  data <= "11111111";  -- 1FA0 = FF
      when "1111110100001" =>  data <= "11111111";  -- 1FA1 = FF
      when "1111110100010" =>  data <= "11111111";  -- 1FA2 = FF
      when "1111110100011" =>  data <= "11111111";  -- 1FA3 = FF
      when "1111110100100" =>  data <= "11111111";  -- 1FA4 = FF
      when "1111110100101" =>  data <= "11111111";  -- 1FA5 = FF
      when "1111110100110" =>  data <= "11111111";  -- 1FA6 = FF
      when "1111110100111" =>  data <= "11111111";  -- 1FA7 = FF
      when "1111110101000" =>  data <= "11111111";  -- 1FA8 = FF
      when "1111110101001" =>  data <= "11111111";  -- 1FA9 = FF
      when "1111110101010" =>  data <= "11111111";  -- 1FAA = FF
      when "1111110101011" =>  data <= "11111111";  -- 1FAB = FF
      when "1111110101100" =>  data <= "11111111";  -- 1FAC = FF
      when "1111110101101" =>  data <= "11111111";  -- 1FAD = FF
      when "1111110101110" =>  data <= "11111111";  -- 1FAE = FF
      when "1111110101111" =>  data <= "11111111";  -- 1FAF = FF
      when "1111110110000" =>  data <= "11111111";  -- 1FB0 = FF
      when "1111110110001" =>  data <= "11111111";  -- 1FB1 = FF
      when "1111110110010" =>  data <= "11111111";  -- 1FB2 = FF
      when "1111110110011" =>  data <= "11111111";  -- 1FB3 = FF
      when "1111110110100" =>  data <= "11111111";  -- 1FB4 = FF
      when "1111110110101" =>  data <= "11111111";  -- 1FB5 = FF
      when "1111110110110" =>  data <= "11111111";  -- 1FB6 = FF
      when "1111110110111" =>  data <= "11111111";  -- 1FB7 = FF
      when "1111110111000" =>  data <= "11111111";  -- 1FB8 = FF
      when "1111110111001" =>  data <= "11111111";  -- 1FB9 = FF
      when "1111110111010" =>  data <= "11111111";  -- 1FBA = FF
      when "1111110111011" =>  data <= "11111111";  -- 1FBB = FF
      when "1111110111100" =>  data <= "11111111";  -- 1FBC = FF
      when "1111110111101" =>  data <= "11111111";  -- 1FBD = FF
      when "1111110111110" =>  data <= "11111111";  -- 1FBE = FF
      when "1111110111111" =>  data <= "11111111";  -- 1FBF = FF
      when "1111111000000" =>  data <= "11111111";  -- 1FC0 = FF
      when "1111111000001" =>  data <= "11111111";  -- 1FC1 = FF
      when "1111111000010" =>  data <= "11111111";  -- 1FC2 = FF
      when "1111111000011" =>  data <= "11111111";  -- 1FC3 = FF
      when "1111111000100" =>  data <= "11111111";  -- 1FC4 = FF
      when "1111111000101" =>  data <= "11111111";  -- 1FC5 = FF
      when "1111111000110" =>  data <= "11111111";  -- 1FC6 = FF
      when "1111111000111" =>  data <= "11111111";  -- 1FC7 = FF
      when "1111111001000" =>  data <= "11111111";  -- 1FC8 = FF
      when "1111111001001" =>  data <= "11111111";  -- 1FC9 = FF
      when "1111111001010" =>  data <= "11111111";  -- 1FCA = FF
      when "1111111001011" =>  data <= "11111111";  -- 1FCB = FF
      when "1111111001100" =>  data <= "11111111";  -- 1FCC = FF
      when "1111111001101" =>  data <= "11111111";  -- 1FCD = FF
      when "1111111001110" =>  data <= "11111111";  -- 1FCE = FF
      when "1111111001111" =>  data <= "11111111";  -- 1FCF = FF
      when "1111111010000" =>  data <= "11111111";  -- 1FD0 = FF
      when "1111111010001" =>  data <= "11111111";  -- 1FD1 = FF
      when "1111111010010" =>  data <= "11111111";  -- 1FD2 = FF
      when "1111111010011" =>  data <= "11111111";  -- 1FD3 = FF
      when "1111111010100" =>  data <= "11111111";  -- 1FD4 = FF
      when "1111111010101" =>  data <= "11111111";  -- 1FD5 = FF
      when "1111111010110" =>  data <= "11111111";  -- 1FD6 = FF
      when "1111111010111" =>  data <= "11111111";  -- 1FD7 = FF
      when "1111111011000" =>  data <= "11111111";  -- 1FD8 = FF
      when "1111111011001" =>  data <= "11111111";  -- 1FD9 = FF
      when "1111111011010" =>  data <= "11111111";  -- 1FDA = FF
      when "1111111011011" =>  data <= "11111111";  -- 1FDB = FF
      when "1111111011100" =>  data <= "11111111";  -- 1FDC = FF
      when "1111111011101" =>  data <= "11111111";  -- 1FDD = FF
      when "1111111011110" =>  data <= "11111111";  -- 1FDE = FF
      when "1111111011111" =>  data <= "11111111";  -- 1FDF = FF
      when "1111111100000" =>  data <= "11111111";  -- 1FE0 = FF
      when "1111111100001" =>  data <= "11111111";  -- 1FE1 = FF
      when "1111111100010" =>  data <= "11111111";  -- 1FE2 = FF
      when "1111111100011" =>  data <= "11111111";  -- 1FE3 = FF
      when "1111111100100" =>  data <= "11111111";  -- 1FE4 = FF
      when "1111111100101" =>  data <= "11111111";  -- 1FE5 = FF
      when "1111111100110" =>  data <= "11111111";  -- 1FE6 = FF
      when "1111111100111" =>  data <= "11111111";  -- 1FE7 = FF
      when "1111111101000" =>  data <= "11111111";  -- 1FE8 = FF
      when "1111111101001" =>  data <= "11111111";  -- 1FE9 = FF
      when "1111111101010" =>  data <= "11111111";  -- 1FEA = FF
      when "1111111101011" =>  data <= "11111111";  -- 1FEB = FF
      when "1111111101100" =>  data <= "11111111";  -- 1FEC = FF
      when "1111111101101" =>  data <= "11111111";  -- 1FED = FF
      when "1111111101110" =>  data <= "11111111";  -- 1FEE = FF
      when "1111111101111" =>  data <= "11111111";  -- 1FEF = FF
      when "1111111110000" =>  data <= "11111111";  -- 1FF0 = FF
      when "1111111110001" =>  data <= "11111111";  -- 1FF1 = FF
      when "1111111110010" =>  data <= "11111111";  -- 1FF2 = FF
      when "1111111110011" =>  data <= "11111111";  -- 1FF3 = FF
      when "1111111110100" =>  data <= "11111111";  -- 1FF4 = FF
      when "1111111110101" =>  data <= "11111111";  -- 1FF5 = FF
      when "1111111110110" =>  data <= "11111111";  -- 1FF6 = FF
      when "1111111110111" =>  data <= "11111111";  -- 1FF7 = FF
      when "1111111111000" =>  data <= "11111111";  -- 1FF8 = FF
      when "1111111111001" =>  data <= "11111111";  -- 1FF9 = FF
      when "1111111111010" =>  data <= "00111000";  -- 1FFA = 38
      when "1111111111011" =>  data <= "11100000";  -- 1FFB = E0
      when "1111111111100" =>  data <= "00000010";  -- 1FFC = 2
      when "1111111111101" =>  data <= "11100000";  -- 1FFD = E0
      when "1111111111110" =>  data <= "00000010";  -- 1FFE = 2
      when "1111111111111" =>  data <= "11100000";  -- 1FFF = E0
      --end_of_rom
      when others =>  data <= "00000000";
    end case;
  end process;

end arch_osrom;

------------------------------------------------------------------------------
------------------------------------------------------------------------------

