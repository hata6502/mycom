is_word(IS_ADD, 0), 	-- 256
is_word(IS_ADD, 0), 	-- 257
is_word(IS_ADD, 0), 	-- 258
is_word(IS_ADD, 0), 	-- 259
is_word(IS_ADD, 0), 	-- 260
is_word(IS_ADD, 0), 	-- 261
is_word(IS_ADD, 0), 	-- 262
is_word(IS_ADD, 0), 	-- 263
is_word(IS_ADD, 0), 	-- 264
is_word(IS_ADD, 0), 	-- 265
is_word(IS_ADD, 0), 	-- 266
is_word(IS_ADD, 0), 	-- 267
is_word(IS_ADD, 0), 	-- 268
is_word(IS_ADD, 0), 	-- 269
is_word(IS_ADD, 0), 	-- 270
is_word(IS_ADD, 0), 	-- 271
is_word(IS_ADD, 0), 	-- 272
is_word(IS_ADD, 0), 	-- 273
is_word(IS_ADD, 0), 	-- 274
is_word(IS_ADD, 0), 	-- 275
is_word(IS_ADD, 0), 	-- 276
is_word(IS_ADD, 0), 	-- 277
is_word(IS_ADD, 0), 	-- 278
is_word(IS_ADD, 0), 	-- 279
is_word(IS_ADD, 0), 	-- 280
is_word(IS_ADD, 0), 	-- 281
is_word(IS_ADD, 0), 	-- 282
is_word(IS_ADD, 0), 	-- 283
is_word(IS_ADD, 0), 	-- 284
is_word(IS_ADD, 0), 	-- 285
is_word(IS_ADD, 0), 	-- 286
is_word(IS_ADD, 0), 	-- 287
is_word(IS_READ, 511), 	-- 288
is_word(IS_WRITE, 2), 	-- 289
is_word(IS_READ, 510), 	-- 290
is_word(IS_WRITE, 2), 	-- 291
is_word(IS_READ, 509), 	-- 292
is_word(IS_WRITE, 2), 	-- 293
is_word(IS_READ, 508), 	-- 294
is_word(IS_WRITE, 507), 	-- 295
is_word(IS_READ, 506), 	-- 296
is_word(IS_WRITE, 2), 	-- 297
is_word(IS_READ, 505), 	-- 298
is_word(IS_WRITE, 2), 	-- 299
is_word(IS_READ, 504), 	-- 300
is_word(IS_WRITE, 2), 	-- 301
is_word(IS_READ, 0), 	-- 302
0, 	-- 303
0, 	-- 304
0, 	-- 305
0, 	-- 306
0, 	-- 307
0, 	-- 308
0, 	-- 309
0, 	-- 310
0, 	-- 311
0, 	-- 312
0, 	-- 313
0, 	-- 314
0, 	-- 315
0, 	-- 316
0, 	-- 317
0, 	-- 318
0, 	-- 319
0, 	-- 320
0, 	-- 321
0, 	-- 322
0, 	-- 323
0, 	-- 324
0, 	-- 325
0, 	-- 326
0, 	-- 327
0, 	-- 328
0, 	-- 329
0, 	-- 330
0, 	-- 331
0, 	-- 332
0, 	-- 333
0, 	-- 334
0, 	-- 335
0, 	-- 336
0, 	-- 337
0, 	-- 338
0, 	-- 339
0, 	-- 340
0, 	-- 341
0, 	-- 342
0, 	-- 343
0, 	-- 344
0, 	-- 345
0, 	-- 346
0, 	-- 347
0, 	-- 348
0, 	-- 349
0, 	-- 350
0, 	-- 351
0, 	-- 352
0, 	-- 353
0, 	-- 354
0, 	-- 355
0, 	-- 356
0, 	-- 357
0, 	-- 358
0, 	-- 359
0, 	-- 360
0, 	-- 361
0, 	-- 362
0, 	-- 363
0, 	-- 364
0, 	-- 365
0, 	-- 366
0, 	-- 367
0, 	-- 368
0, 	-- 369
0, 	-- 370
0, 	-- 371
0, 	-- 372
0, 	-- 373
0, 	-- 374
0, 	-- 375
0, 	-- 376
0, 	-- 377
0, 	-- 378
0, 	-- 379
0, 	-- 380
0, 	-- 381
0, 	-- 382
0, 	-- 383
0, 	-- 384
0, 	-- 385
0, 	-- 386
0, 	-- 387
0, 	-- 388
0, 	-- 389
0, 	-- 390
0, 	-- 391
0, 	-- 392
0, 	-- 393
0, 	-- 394
0, 	-- 395
0, 	-- 396
0, 	-- 397
0, 	-- 398
0, 	-- 399
0, 	-- 400
0, 	-- 401
0, 	-- 402
0, 	-- 403
0, 	-- 404
0, 	-- 405
0, 	-- 406
0, 	-- 407
0, 	-- 408
0, 	-- 409
0, 	-- 410
0, 	-- 411
0, 	-- 412
0, 	-- 413
0, 	-- 414
0, 	-- 415
0, 	-- 416
0, 	-- 417
0, 	-- 418
0, 	-- 419
0, 	-- 420
0, 	-- 421
0, 	-- 422
0, 	-- 423
0, 	-- 424
0, 	-- 425
0, 	-- 426
0, 	-- 427
0, 	-- 428
0, 	-- 429
0, 	-- 430
0, 	-- 431
0, 	-- 432
0, 	-- 433
0, 	-- 434
0, 	-- 435
0, 	-- 436
0, 	-- 437
0, 	-- 438
0, 	-- 439
0, 	-- 440
0, 	-- 441
0, 	-- 442
0, 	-- 443
0, 	-- 444
0, 	-- 445
0, 	-- 446
0, 	-- 447
0, 	-- 448
0, 	-- 449
0, 	-- 450
0, 	-- 451
0, 	-- 452
0, 	-- 453
0, 	-- 454
0, 	-- 455
0, 	-- 456
0, 	-- 457
0, 	-- 458
0, 	-- 459
0, 	-- 460
0, 	-- 461
0, 	-- 462
0, 	-- 463
0, 	-- 464
0, 	-- 465
0, 	-- 466
0, 	-- 467
0, 	-- 468
0, 	-- 469
0, 	-- 470
0, 	-- 471
0, 	-- 472
0, 	-- 473
0, 	-- 474
0, 	-- 475
0, 	-- 476
0, 	-- 477
0, 	-- 478
0, 	-- 479
0, 	-- 480
0, 	-- 481
0, 	-- 482
0, 	-- 483
0, 	-- 484
0, 	-- 485
0, 	-- 486
0, 	-- 487
0, 	-- 488
0, 	-- 489
0, 	-- 490
0, 	-- 491
0, 	-- 492
0, 	-- 493
0, 	-- 494
0, 	-- 495
0, 	-- 496
0, 	-- 497
0, 	-- 498
0, 	-- 499
0, 	-- 500
0, 	-- 501
0, 	-- 502
0, 	-- 503
0, 	-- 504
1280, 	-- 505
0, 	-- 506
0, 	-- 507
0, 	-- 508
0, 	-- 509
1024, 	-- 510
296	-- 511
