LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

ENTITY crom IS
	PORT (
		chr : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		row : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		col : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		dot : OUT STD_LOGIC
	);
END crom;
ARCHITECTURE Behavioral OF crom IS

	SUBTYPE crom_row IS STD_LOGIC_VECTOR(0 TO 7);
	TYPE crom_chr IS ARRAY (0 TO 7) OF crom_row;
	TYPE crom IS ARRAY (0 TO 255) OF crom_chr;
	CONSTANT crom_1 : crom :=
	(
	(
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (-- SP
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (-- !
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00000000",
	"00010000",
	"00000000"
	), (-- "
	"11011000",
	"01001000",
	"10010000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (-- #
	"00010100",
	"01111110",
	"00101000",
	"00101000",
	"00101000",
	"11111100",
	"01010000",
	"00000000"
	), (-- $
	"00001000",
	"00111110",
	"01001000",
	"00111100",
	"00010010",
	"01111100",
	"00010000",
	"00000000"
	), (-- %
	"01000010",
	"10100100",
	"01001000",
	"00010000",
	"00100100",
	"01001010",
	"10000100",
	"00000000"
	), (-- &
	"00110000",
	"01001000",
	"01010000",
	"00100100",
	"01010100",
	"10001000",
	"01110110",
	"00000000"
	), (-- '
	"11000000",
	"01000000",
	"10000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (-- (
	"00000010",
	"00000100",
	"00001000",
	"00001000",
	"00001000",
	"00000100",
	"00000010",
	"00000000"
	), (-- )
	"10000000",
	"01000000",
	"00100000",
	"00100000",
	"00100000",
	"01000000",
	"10000000",
	"00000000"
	), (-- *
	"00010000",
	"01010100",
	"00111000",
	"00010000",
	"00111000",
	"01010100",
	"00010000",
	"00000000"
	), (-- +
	"00010000",
	"00010000",
	"00010000",
	"11111110",
	"00010000",
	"00010000",
	"00010000",
	"00000000"
	), (-- ,
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11000000",
	"01000000",
	"10000000",
	"00000000"
	), (-- -
	"00000000",
	"00000000",
	"00000000",
	"11111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (-- .
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11000000",
	"11000000",
	"00000000"
	), (-- /
	"00000010",
	"00000100",
	"00001000",
	"00010000",
	"00100000",
	"01000000",
	"10000000",
	"00000000"
	), (-- 0
	"00111100",
	"01000010",
	"01000010",
	"01000010",
	"01000010",
	"01000010",
	"00111100",
	"00000000"
	), (
	"00010000",
	"00110000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00111000",
	"00000000"
	), (
	"00111100",
	"01000010",
	"00000010",
	"00001100",
	"00110000",
	"01000000",
	"01111110",
	"00000000"
	), (
	"00111100",
	"01000010",
	"00000010",
	"00011100",
	"00000010",
	"01000010",
	"00111100",
	"00000000"
	), (
	"00000100",
	"00001100",
	"00010100",
	"00100100",
	"01000100",
	"01111110",
	"00000100",
	"00000000"
	), (
	"01111110",
	"01000000",
	"01111100",
	"01000010",
	"00000010",
	"01000010",
	"00111100",
	"00000000"
	), (
	"00111100",
	"01000010",
	"01000000",
	"01111100",
	"01000010",
	"01000010",
	"00111100",
	"00000000"
	), (
	"01111110",
	"00000010",
	"00000100",
	"00001000",
	"00001000",
	"00010000",
	"00010000",
	"00000000"
	), (
	"00111100",
	"01000010",
	"01000010",
	"00111100",
	"01000010",
	"01000010",
	"00111100",
	"00000000"
	), (-- 9
	"00111100",
	"01000010",
	"01000010",
	"00111110",
	"00000010",
	"01000010",
	"00111100",
	"00000000"
	), (-- :
	"00000000",
	"00110000",
	"00110000",
	"00000000",
	"00110000",
	"00110000",
	"00000000",
	"00000000"
	), (-- ;
	"00000000",
	"00110000",
	"00110000",
	"00000000",
	"00110000",
	"00010000",
	"00100000",
	"00000000"
	), (-- <
	"00000010",
	"00000100",
	"00001000",
	"00010000",
	"00001000",
	"00000100",
	"00000010",
	"00000000"
	), (-- =
	"00000000",
	"00000000",
	"11111110",
	"00000000",
	"11111110",
	"00000000",
	"00000000",
	"00000000"
	), (-- >
	"10000000",
	"01000000",
	"00100000",
	"00010000",
	"00100000",
	"01000000",
	"10000000",
	"00000000"
	), (-- ?
	"00111100",
	"01000010",
	"00000010",
	"00001100",
	"00010000",
	"00000000",
	"00010000",
	"00000000"
	), (-- @
	"00111000",
	"01000100",
	"10011010",
	"10101010",
	"10110100",
	"01000000",
	"00111000",
	"00000000"
	), (-- A
	"00010000",
	"00101000",
	"00101000",
	"01000100",
	"01111100",
	"10000010",
	"10000010",
	"00000000"
	), (
	"01111100",
	"01000010",
	"01000010",
	"01111100",
	"01000010",
	"01000010",
	"01111100",
	"00000000"
	), (
	"00011100",
	"00100010",
	"01000000",
	"01000000",
	"01000000",
	"00100010",
	"00011100",
	"00000000"
	), (
	"01111000",
	"01000100",
	"01000010",
	"01000010",
	"01000010",
	"01000100",
	"01111000",
	"00000000"
	), (
	"01111110",
	"01000000",
	"01000000",
	"01111100",
	"01000000",
	"01000000",
	"01111110",
	"00000000"
	), (
	"01111110",
	"01000000",
	"01000000",
	"01111100",
	"01000000",
	"01000000",
	"01000000",
	"00000000"
	), (
	"00011100",
	"00100010",
	"01000000",
	"01001110",
	"01000010",
	"00100010",
	"00011100",
	"00000000"
	), (
	"01000010",
	"01000010",
	"01000010",
	"01111110",
	"01000010",
	"01000010",
	"01000010",
	"00000000"
	), (
	"00111000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00111000",
	"00000000"
	), (
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"01000010",
	"00111100",
	"00000000"
	), (
	"01000010",
	"01000100",
	"01001000",
	"01010000",
	"01101000",
	"01000100",
	"01000010",
	"00000000"
	), (
	"01000000",
	"01000000",
	"01000000",
	"01000000",
	"01000000",
	"01000000",
	"01111110",
	"00000000"
	), (
	"10000010",
	"11000110",
	"10101010",
	"10101010",
	"10010010",
	"10010010",
	"10000010",
	"00000000"
	), (
	"01000010",
	"01100010",
	"01010010",
	"01001010",
	"01000110",
	"01000010",
	"01000010",
	"00000000"
	), (
	"00011000",
	"00100100",
	"01000010",
	"01000010",
	"01000010",
	"00100100",
	"00011000",
	"00000000"
	), (
	"01111100",
	"01000010",
	"01000010",
	"01111100",
	"01000000",
	"01000000",
	"01000000",
	"00000000"
	), (
	"00011000",
	"00100100",
	"01000010",
	"01000010",
	"01001010",
	"00100100",
	"00011010",
	"00000000"
	), (
	"01111100",
	"01000010",
	"01000010",
	"01111100",
	"01001000",
	"01000100",
	"01000010",
	"00000000"
	), (
	"00111100",
	"01000010",
	"01000000",
	"00111100",
	"00000010",
	"01000010",
	"00111100",
	"00000000"
	), (
	"11111110",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00000000"
	), (
	"01000010",
	"01000010",
	"01000010",
	"01000010",
	"01000010",
	"01000010",
	"00111100",
	"00000000"
	), (
	"10000010",
	"10000010",
	"01000100",
	"01000100",
	"00101000",
	"00101000",
	"00010000",
	"00000000"
	), (
	"10000010",
	"10010010",
	"10010010",
	"10101010",
	"10101010",
	"01000100",
	"01000100",
	"00000000"
	), (
	"10000010",
	"01000100",
	"00101000",
	"00010000",
	"00101000",
	"01000100",
	"10000010",
	"00000000"
	), (
	"10000010",
	"01000100",
	"00101000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00000000"
	), (-- Z
	"01111110",
	"00000010",
	"00000100",
	"00001000",
	"00010000",
	"00100000",
	"01111110",
	"00000000"
	), (-- [
	"00001110",
	"00001000",
	"00001000",
	"00001000",
	"00001000",
	"00001000",
	"00001110",
	"00000000"
	), (-- \
	"10000000",
	"01000000",
	"00100000",
	"00010000",
	"00001000",
	"00000100",
	"00000010",
	"00000000"
	), (-- ]
	"11100000",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"11100000",
	"00000000"
	), (-- ^
	"00010000",
	"00101000",
	"01000100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (-- _
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111110",
	"00000000"
	), (-- `
	"10000000",
	"01000000",
	"00100000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (-- a
	"00000000",
	"00000000",
	"00111000",
	"00000100",
	"00111100",
	"01000100",
	"00111100",
	"00000000"
	), (
	"01000000",
	"01000000",
	"01011000",
	"01100100",
	"01000100",
	"01000100",
	"01111000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00111000",
	"01000100",
	"01000000",
	"01000100",
	"00111000",
	"00000000"
	), (
	"00000100",
	"00000100",
	"00110100",
	"01001100",
	"01000100",
	"01000100",
	"00111100",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00111000",
	"01000100",
	"01111100",
	"01000000",
	"00111000",
	"00000000"
	), (
	"00001100",
	"00010000",
	"00111000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00111100",
	"01000100",
	"00111100",
	"00000100",
	"00111000",
	"00000000"
	), (
	"01000000",
	"01000000",
	"01011000",
	"01100100",
	"01000100",
	"01000100",
	"01000100",
	"00000000"
	), (
	"00010000",
	"00000000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00000000"
	), (
	"00001000",
	"00000000",
	"00001000",
	"00001000",
	"00001000",
	"01001000",
	"00110000",
	"00000000"
	), (
	"00100000",
	"00100000",
	"00100100",
	"00101000",
	"00110000",
	"00101000",
	"00100100",
	"00000000"
	), (
	"00110000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"01101000",
	"01010100",
	"01010100",
	"01010100",
	"01010100",
	"00000000"
	), (
	"00000000",
	"00000000",
	"01011000",
	"01100100",
	"01000100",
	"01000100",
	"01000100",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00111000",
	"01000100",
	"01000100",
	"01000100",
	"00111000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"01111000",
	"01000100",
	"01111000",
	"01000000",
	"01000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00111100",
	"01000100",
	"00111100",
	"00000100",
	"00000100",
	"00000000"
	), (
	"00000000",
	"00000000",
	"01011000",
	"01100100",
	"01000000",
	"01000000",
	"01000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00111100",
	"01000000",
	"00111000",
	"00000100",
	"01111000",
	"00000000"
	), (
	"00000000",
	"00100000",
	"01111000",
	"00100000",
	"00100000",
	"00100100",
	"00011000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"01000100",
	"01000100",
	"01000100",
	"01001100",
	"00110100",
	"00000000"
	), (
	"00000000",
	"00000000",
	"01000100",
	"01000100",
	"00101000",
	"00101000",
	"00010000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"01000100",
	"01010100",
	"01010100",
	"00101000",
	"00101000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"01000100",
	"00101000",
	"00010000",
	"00101000",
	"01000100",
	"00000000"
	), (
	"00000000",
	"00000000",
	"01000100",
	"00101000",
	"00101000",
	"00010000",
	"01100000",
	"00000000"
	), (-- z
	"00000000",
	"00000000",
	"01111100",
	"00001000",
	"00010000",
	"00100000",
	"01111100",
	"00000000"
	), (-- {
	"00000110",
	"00001000",
	"00001000",
	"00010000",
	"00001000",
	"00001000",
	"00000110",
	"00000000"
	), (-- |
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00000000"
	), (-- }
	"11000000",
	"00100000",
	"00100000",
	"00010000",
	"00100000",
	"00100000",
	"11000000",
	"00000000"
	), (-- ~
	"00000000",
	"00000000",
	"01100000",
	"10010010",
	"00001100",
	"00000000",
	"00000000",
	"00000000"
	), (-- DEL
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	),

	(
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	),

	(-- SP
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (-- �
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01000000",
	"10100000",
	"01000000",
	"00000000"
	), (-- �
	"00011110",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00000000",
	"00000000"
	), (-- �
	"00000000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"11110000",
	"00000000"
	), (-- �
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"10000000",
	"01000000",
	"00000000"
	), (-- �
	"00000000",
	"00000000",
	"00000000",
	"00110000",
	"00110000",
	"00000000",
	"00000000",
	"00000000"
	), (-- ��
	"01111110",
	"00000010",
	"00111110",
	"00000010",
	"00000100",
	"00001000",
	"00110000",
	"00000000"
	), (-- �@
	"00000000",
	"00000000",
	"01111100",
	"00010100",
	"00011000",
	"00010000",
	"00100000",
	"00000000"
	), (-- �B
	"00000000",
	"00000000",
	"00000100",
	"00001000",
	"00011000",
	"01101000",
	"00001000",
	"00000000"
	), (-- �D
	"00000000",
	"00000000",
	"00010000",
	"01111100",
	"01000100",
	"00001000",
	"00110000",
	"00000000"
	), (-- �F
	"00000000",
	"00000000",
	"00000000",
	"00111000",
	"00010000",
	"00010000",
	"01111100",
	"00000000"
	), (-- �H
	"00000000",
	"00000000",
	"00001000",
	"01111100",
	"00011000",
	"01101000",
	"00011000",
	"00000000"
	), (-- ��
	"00000000",
	"00000000",
	"00100000",
	"00111100",
	"01100100",
	"00010000",
	"00010000",
	"00000000"
	), (-- ��
	"00000000",
	"00000000",
	"00000000",
	"00111000",
	"00001000",
	"00001000",
	"01111100",
	"00000000"
	), (-- ��
	"00000000",
	"00000000",
	"00111100",
	"00000100",
	"00011100",
	"00000100",
	"00111100",
	"00000000"
	), (-- �b
	"00000000",
	"00000000",
	"00000000",
	"01010100",
	"01010100",
	"00001000",
	"00110000",
	"00000000"
	), (-- �
	"00000000",
	"00000000",
	"10000000",
	"01111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (-- �A
	"01111110",
	"00000010",
	"00010100",
	"00011000",
	"00010000",
	"00010000",
	"00100000",
	"00000000"
	), (-- �C
	"00000010",
	"00000100",
	"00001000",
	"00011000",
	"01101000",
	"00001000",
	"00001000",
	"00000000"
	), (-- �E
	"00010000",
	"01111110",
	"01000010",
	"00000010",
	"00000100",
	"00001000",
	"00110000",
	"00000000"
	), (-- �G
	"00000000",
	"01111100",
	"00010000",
	"00010000",
	"00010000",
	"11111110",
	"00000000",
	"00000000"
	), (-- �I
	"00001000",
	"11111110",
	"00001000",
	"00011000",
	"00101000",
	"11001000",
	"00011000",
	"00000000"
	), (-- �J
	"00010000",
	"01111110",
	"00010010",
	"00010010",
	"00010010",
	"00100010",
	"01000110",
	"00000000"
	), (-- �L
	"00010000",
	"01111100",
	"00010000",
	"00010000",
	"01111110",
	"00001000",
	"00001000",
	"00000000"
	), (-- �N
	"00010000",
	"00011110",
	"00100010",
	"01000010",
	"00000100",
	"00001000",
	"00110000",
	"00000000"
	), (-- �P
	"01000000",
	"01111110",
	"01001000",
	"10001000",
	"00001000",
	"00010000",
	"00100000",
	"00000000"
	), (-- �R
	"00000000",
	"01111110",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"01111110",
	"00000000"
	), (-- �T
	"00100100",
	"11111110",
	"00100100",
	"00100100",
	"00000100",
	"00001000",
	"00110000",
	"00000000"
	), (-- �V
	"01000000",
	"00100000",
	"01000010",
	"00100010",
	"00000100",
	"00001000",
	"01110000",
	"00000000"
	), (-- �X
	"00000000",
	"01111100",
	"00000100",
	"00001000",
	"00001000",
	"00110100",
	"11000010",
	"00000000"
	), (-- �Z
	"00100000",
	"00100000",
	"11111110",
	"00100010",
	"00100100",
	"00100000",
	"00011110",
	"00000000"
	), (-- �\
	"01000010",
	"00100010",
	"00100010",
	"00000010",
	"00000100",
	"00001000",
	"00110000",
	"00000000"
	), (-- �^
	"00010000",
	"00011110",
	"00100010",
	"01011010",
	"00000100",
	"00001000",
	"00110000",
	"00000000"
	), (-- �`
	"00001100",
	"01110000",
	"00010000",
	"11111110",
	"00010000",
	"00010000",
	"00100000",
	"00000000"
	), (-- �
	"00000000",
	"10100010",
	"01010010",
	"01010010",
	"00000100",
	"00001000",
	"00110000",
	"00000000"
	), (-- �e
	"01111100",
	"00000000",
	"11111110",
	"00010000",
	"00010000",
	"00010000",
	"00100000",
	"00000000"
	), (-- �g
	"00100000",
	"00100000",
	"00100000",
	"00111000",
	"00100100",
	"00100000",
	"00100000",
	"00000000"
	), (-- �i
	"00010000",
	"00010000",
	"11111110",
	"00010000",
	"00010000",
	"00100000",
	"01000000",
	"00000000"
	), (-- �j
	"00000000",
	"01111100",
	"00000000",
	"00000000",
	"00000000",
	"11111110",
	"00000000",
	"00000000"
	), (-- �k
	"01111100",
	"00000100",
	"00110100",
	"00001000",
	"00011000",
	"00100100",
	"11000000",
	"00000000"
	), (-- �l
	"00010000",
	"01111100",
	"00001000",
	"00010000",
	"00110100",
	"11010010",
	"00010000",
	"00000000"
	), (-- �m
	"00000100",
	"00000100",
	"00000100",
	"00001000",
	"00010000",
	"00100000",
	"11000000",
	"00000000"
	), (-- �n
	"00000000",
	"00101000",
	"00100100",
	"00100100",
	"01000010",
	"01000010",
	"10000010",
	"00000000"
	), (-- �q
	"01000000",
	"01000000",
	"01000110",
	"01111000",
	"01000000",
	"01000000",
	"00111110",
	"00000000"
	), (-- �t
	"00000000",
	"01111110",
	"00000010",
	"00000010",
	"00000100",
	"00001000",
	"00110000",
	"00000000"
	), (-- �w
	"00000000",
	"00100000",
	"01010000",
	"10001000",
	"00000100",
	"00000010",
	"00000000",
	"00000000"
	), (-- �z
	"00010000",
	"00010000",
	"11111110",
	"00010000",
	"01010100",
	"10010010",
	"00110000",
	"00000000"
	), (-- �}
	"00000000",
	"11111110",
	"00000010",
	"00000100",
	"00101000",
	"00010000",
	"00001000",
	"00000000"
	), (-- �~
	"01110000",
	"00001100",
	"00100000",
	"00011000",
	"00000000",
	"01110000",
	"00001100",
	"00000000"
	), (-- ��
	"00010000",
	"00010000",
	"00100000",
	"00100000",
	"01001000",
	"01000100",
	"11111010",
	"00000000"
	), (-- ��
	"00000100",
	"00000100",
	"01110100",
	"00001000",
	"00010100",
	"00100100",
	"11000000",
	"00000000"
	), (-- ��
	"00111100",
	"00010000",
	"00010000",
	"01111110",
	"00010000",
	"00010000",
	"00001110",
	"00000000"
	), (-- ��
	"00100000",
	"00101110",
	"11110010",
	"00100100",
	"00010000",
	"00010000",
	"00010000",
	"00000000"
	), (-- ��
	"00000000",
	"01111000",
	"00001000",
	"00001000",
	"00001000",
	"11111110",
	"00000000",
	"00000000"
	), (-- ��
	"00000000",
	"01111110",
	"00000010",
	"00111110",
	"00000010",
	"00000010",
	"01111110",
	"00000000"
	), (-- ��
	"00111100",
	"00000000",
	"01111110",
	"00000010",
	"00000100",
	"00001000",
	"00110000",
	"00000000"
	), (-- ��
	"01000100",
	"01000100",
	"01000100",
	"01000100",
	"00000100",
	"00001000",
	"00110000",
	"00000000"
	), (-- ��
	"00001000",
	"00101000",
	"00101000",
	"00101000",
	"00101010",
	"01001100",
	"10001000",
	"00000000"
	), (-- ��
	"00100000",
	"00100000",
	"00100000",
	"00100010",
	"00100100",
	"00101000",
	"00110000",
	"00000000"
	), (-- ��
	"00000000",
	"01111110",
	"01000010",
	"01000010",
	"01000010",
	"01000010",
	"01111110",
	"00000000"
	), (-- ��
	"00000000",
	"01111110",
	"01000010",
	"00000010",
	"00000100",
	"00001000",
	"00110000",
	"00000000"
	), (-- ��
	"01000000",
	"00100000",
	"00000010",
	"00000010",
	"00000100",
	"00001000",
	"01110000",
	"00000000"
	), (-- �
	"10100000",
	"01010000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (-- �
	"01000000",
	"10100000",
	"01000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	),

	(
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	), (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000"
	)

	);

BEGIN
	dot <= crom_1(conv_integer(chr))(conv_integer(row))(conv_integer(col));
END Behavioral;