iconv input.asm -f utf8 -t sjis > input.c
gcc -E -P input.c > input_pre.asm
rm input.c
./asm < input_pre.asm
is_word(IS_ADD, 3), 	-- 256
is_word(IS_ADD, 3), 	-- 257
is_word(IS_ADD, 3), 	-- 258
is_word(IS_ADD, 3), 	-- 259
is_word(IS_ADD, 3), 	-- 260
is_word(IS_ADD, 3), 	-- 261
is_word(IS_ADD, 3), 	-- 262
is_word(IS_ADD, 3), 	-- 263
is_word(IS_ADD, 3), 	-- 264
is_word(IS_ADD, 3), 	-- 265
is_word(IS_ADD, 3), 	-- 266
is_word(IS_ADD, 3), 	-- 267
is_word(IS_ADD, 3), 	-- 268
is_word(IS_ADD, 3), 	-- 269
is_word(IS_ADD, 3), 	-- 270
is_word(IS_ADD, 3), 	-- 271
is_word(IS_ADD, 3), 	-- 272
is_word(IS_ADD, 3), 	-- 273
is_word(IS_ADD, 3), 	-- 274
is_word(IS_ADD, 3), 	-- 275
is_word(IS_ADD, 3), 	-- 276
is_word(IS_ADD, 3), 	-- 277
is_word(IS_ADD, 3), 	-- 278
is_word(IS_ADD, 3), 	-- 279
is_word(IS_ADD, 3), 	-- 280
is_word(IS_ADD, 3), 	-- 281
is_word(IS_ADD, 3), 	-- 282
is_word(IS_ADD, 3), 	-- 283
is_word(IS_ADD, 3), 	-- 284
is_word(IS_ADD, 3), 	-- 285
is_word(IS_ADD, 3), 	-- 286
is_word(IS_ADD, 3), 	-- 287
is_word(IS_READ, 767), 	-- 288
is_word(IS_WRITE, 766), 	-- 289
is_word(IS_READ, 66), 	-- 290
is_word(IS_READ, 108), 	-- 291
is_word(IS_READ, 117), 	-- 292
is_word(IS_READ, 101), 	-- 293
is_word(IS_READ, 72), 	-- 294
is_word(IS_READ, 111), 	-- 295
is_word(IS_READ, 111), 	-- 296
is_word(IS_READ, 100), 	-- 297
is_word(IS_READ, 32), 	-- 298
is_word(IS_READ, 67), 	-- 299
is_word(IS_READ, 111), 	-- 300
is_word(IS_READ, 109), 	-- 301
is_word(IS_READ, 112), 	-- 302
is_word(IS_READ, 117), 	-- 303
is_word(IS_READ, 116), 	-- 304
is_word(IS_READ, 101), 	-- 305
is_word(IS_READ, 114), 	-- 306
is_word(IS_READ, 32), 	-- 307
is_word(IS_READ, 32), 	-- 308
is_word(IS_READ, 210), 	-- 309
is_word(IS_READ, 178), 	-- 310
is_word(IS_READ, 219), 	-- 311
is_word(IS_READ, 32), 	-- 312
is_word(IS_READ, 190), 	-- 313
is_word(IS_READ, 178), 	-- 314
is_word(IS_READ, 190), 	-- 315
is_word(IS_READ, 178), 	-- 316
is_word(IS_READ, 32), 	-- 317
is_word(IS_READ, 204), 	-- 318
is_word(IS_READ, 223), 	-- 319
is_word(IS_READ, 219), 	-- 320
is_word(IS_READ, 184), 	-- 321
is_word(IS_READ, 222), 	-- 322
is_word(IS_READ, 215), 	-- 323
is_word(IS_READ, 209), 	-- 324
is_word(IS_READ, 0), 	-- 325
is_word(IS_READ, 206), 	-- 326
is_word(IS_READ, 222), 	-- 327
is_word(IS_READ, 192), 	-- 328
is_word(IS_READ, 221), 	-- 329
is_word(IS_READ, 166), 	-- 330
is_word(IS_READ, 32), 	-- 331
is_word(IS_READ, 181), 	-- 332
is_word(IS_READ, 190), 	-- 333
is_word(IS_READ, 33), 	-- 334
is_word(IS_READ, 32), 	-- 335
is_word(IS_READ, 0), 	-- 336
is_word(IS_READ, 219), 	-- 337
is_word(IS_READ, 0), 	-- 338
is_word(IS_READ, 765), 	-- 339
is_word(IS_WRITE, 2), 	-- 340
is_word(IS_READ, 764), 	-- 341
is_word(IS_WRITE, 2), 	-- 342
is_word(IS_READ, 763), 	-- 343
is_word(IS_WRITE, 2), 	-- 344
is_word(IS_READ, 762), 	-- 345
is_word(IS_WRITE, 761), 	-- 346
is_word(IS_READ, 760), 	-- 347
is_word(IS_WRITE, 2), 	-- 348
is_word(IS_READ, 759), 	-- 349
is_word(IS_WRITE, 2), 	-- 350
is_word(IS_READ, 758), 	-- 351
is_word(IS_WRITE, 2), 	-- 352
is_word(IS_READ, 757), 	-- 353
is_word(IS_WRITE, 756), 	-- 354
is_word(IS_READ, 7), 	-- 355
is_word(IS_EQ, 755), 	-- 356
is_word(IS_BRANCH, 754), 	-- 357
is_word(IS_READ, 753), 	-- 358
is_word(IS_WRITE, 752), 	-- 359
is_word(IS_READ, 196), 	-- 360
is_word(IS_GTE, 751), 	-- 361
is_word(IS_BRANCH, 750), 	-- 362
is_word(IS_READ, 749), 	-- 363
is_word(IS_WRITE, 748), 	-- 364
is_word(IS_READ, 197), 	-- 365
is_word(IS_GTE, 747), 	-- 366
is_word(IS_BRANCH, 746), 	-- 367
is_word(IS_READ, 196), 	-- 368
is_word(IS_EQ, 745), 	-- 369
is_word(IS_BRANCH, 744), 	-- 370
is_word(IS_READ, 196), 	-- 371
is_word(IS_EQ, 743), 	-- 372
is_word(IS_BRANCH, 742), 	-- 373
is_word(IS_READ, 197), 	-- 374
is_word(IS_EQ, 741), 	-- 375
is_word(IS_BRANCH, 740), 	-- 376
is_word(IS_READ, 197), 	-- 377
is_word(IS_EQ, 739), 	-- 378
is_word(IS_BRANCH, 738), 	-- 379
is_word(IS_READ, 196), 	-- 380
is_word(IS_OR, 197), 	-- 381
is_word(IS_AND, 737), 	-- 382
is_word(IS_EQ, 736), 	-- 383
is_word(IS_BRANCH, 735), 	-- 384
is_word(IS_READ, 734), 	-- 385
is_word(IS_WRITE, 733), 	-- 386
is_word(IS_READ, 196), 	-- 387
is_word(IS_MUL, 732), 	-- 388
is_word(IS_ADD, 197), 	-- 389
is_word(IS_ADD, 731), 	-- 390
is_word(IS_WRITE, 730), 	-- 391
is_word(IS_READ, 729), 	-- 392
is_word(IS_WRITE, 2), 	-- 393
is_word(IS_READ, 192), 	-- 394
is_word(IS_WRITE, 2), 	-- 395
is_word(IS_READ, 728), 	-- 396
is_word(IS_WRITE, 2), 	-- 397
is_word(IS_READ, 727), 	-- 398
is_word(IS_WRITE, 726), 	-- 399
is_word(IS_READ, 197), 	-- 400
is_word(IS_ADD, 725), 	-- 401
is_word(IS_WRITE, 724), 	-- 402
is_word(IS_READ, 723), 	-- 403
is_word(IS_WRITE, 722), 	-- 404
is_word(IS_READ, 196), 	-- 405
is_word(IS_ADD, 721), 	-- 406
is_word(IS_WRITE, 720), 	-- 407
is_word(IS_READ, 719), 	-- 408
is_word(IS_WRITE, 718), 	-- 409
is_word(IS_READ, 717), 	-- 410
is_word(IS_WRITE, 716), 	-- 411
is_word(IS_READ, 196), 	-- 412
is_word(IS_GTE, 715), 	-- 413
is_word(IS_BRANCH, 714), 	-- 414
is_word(IS_READ, 3), 	-- 415
is_word(IS_AND, 713), 	-- 416
is_word(IS_WRITE, 712), 	-- 417
is_word(IS_READ, 711), 	-- 418
is_word(IS_WRITE, 2), 	-- 419
is_word(IS_READ, 197), 	-- 420
is_word(IS_WRITE, 2), 	-- 421
is_word(IS_READ, 710), 	-- 422
is_word(IS_WRITE, 2), 	-- 423
is_word(IS_READ, 196), 	-- 424
is_word(IS_WRITE, 2), 	-- 425
is_word(IS_READ, 709), 	-- 426
is_word(IS_WRITE, 708), 	-- 427
is_word(IS_READ, 248), 	-- 428
is_word(IS_BRANCH, 707), 	-- 429
is_word(IS_READ, 196), 	-- 430
is_word(IS_ADD, 706), 	-- 431
is_word(IS_WRITE, 705), 	-- 432
is_word(IS_READ, 704), 	-- 433
is_word(IS_WRITE, 703), 	-- 434
is_word(IS_READ, 702), 	-- 435
is_word(IS_WRITE, 701), 	-- 436
is_word(IS_READ, 196), 	-- 437
is_word(IS_GTE, 700), 	-- 438
is_word(IS_BRANCH, 699), 	-- 439
is_word(IS_READ, 698), 	-- 440
is_word(IS_WRITE, 697), 	-- 441
is_word(IS_READ, 197), 	-- 442
is_word(IS_GTE, 696), 	-- 443
is_word(IS_BRANCH, 695), 	-- 444
is_word(IS_READ, 3), 	-- 445
is_word(IS_AND, 694), 	-- 446
is_word(IS_WRITE, 693), 	-- 447
is_word(IS_EQ, 692), 	-- 448
is_word(IS_BRANCH, 691), 	-- 449
is_word(IS_READ, 690), 	-- 450
is_word(IS_WRITE, 2), 	-- 451
is_word(IS_READ, 192), 	-- 452
is_word(IS_WRITE, 2), 	-- 453
is_word(IS_READ, 196), 	-- 454
is_word(IS_WRITE, 2), 	-- 455
is_word(IS_READ, 197), 	-- 456
is_word(IS_WRITE, 2), 	-- 457
is_word(IS_READ, 689), 	-- 458
is_word(IS_WRITE, 688), 	-- 459
is_word(IS_READ, 248), 	-- 460
is_word(IS_BRANCH, 687), 	-- 461
is_word(IS_READ, 197), 	-- 462
is_word(IS_ADD, 686), 	-- 463
is_word(IS_WRITE, 685), 	-- 464
is_word(IS_READ, 684), 	-- 465
is_word(IS_WRITE, 683), 	-- 466
is_word(IS_READ, 196), 	-- 467
is_word(IS_ADD, 682), 	-- 468
is_word(IS_WRITE, 681), 	-- 469
is_word(IS_READ, 680), 	-- 470
is_word(IS_WRITE, 679), 	-- 471
is_word(IS_READ, 7), 	-- 472
is_word(IS_DIV, 678), 	-- 473
is_word(IS_ADD, 677), 	-- 474
is_word(IS_WRITE, 676), 	-- 475
is_word(IS_READ, 7), 	-- 476
is_word(IS_AND, 675), 	-- 477
is_word(IS_ADD, 674), 	-- 478
is_word(IS_WRITE, 673), 	-- 479
is_word(IS_READ, 672), 	-- 480
is_word(IS_WRITE, 671), 	-- 481
is_word(IS_READ, 2), 	-- 482
is_word(IS_WRITE, 670), 	-- 483
is_word(IS_ADD, 3), 	-- 484
is_word(IS_WRITE, 669), 	-- 485
is_word(IS_READ, 2), 	-- 486
is_word(IS_WRITE, 668), 	-- 487
is_word(IS_ADD, 3), 	-- 488
is_word(IS_WRITE, 667), 	-- 489
is_word(IS_READ, 2), 	-- 490
is_word(IS_WRITE, 666), 	-- 491
is_word(IS_ADD, 3), 	-- 492
is_word(IS_WRITE, 665), 	-- 493
is_word(IS_READ, 251), 	-- 494
is_word(IS_MUL, 664), 	-- 495
is_word(IS_ADD, 250), 	-- 496
is_word(IS_ADD, 663), 	-- 497
is_word(IS_WRITE, 662), 	-- 498
is_word(IS_READ, 252), 	-- 499
is_word(IS_NEQ, 661), 	-- 500
is_word(IS_BRANCH, 660), 	-- 501
is_word(IS_READ, 249), 	-- 502
is_word(IS_SUB, 659), 	-- 503
is_word(IS_WRITE, 658), 	-- 504
is_word(IS_READ, 657), 	-- 505
is_word(IS_WRITE, 656), 	-- 506
is_word(IS_READ, 252), 	-- 507
is_word(IS_NEQ, 655), 	-- 508
is_word(IS_BRANCH, 654), 	-- 509
is_word(IS_READ, 249), 	-- 510
is_word(IS_ADD, 653), 	-- 511
is_word(IS_WRITE, 652), 	-- 512
is_word(IS_READ, 651), 	-- 513
is_word(IS_WRITE, 650), 	-- 514
is_word(IS_READ, 252), 	-- 515
is_word(IS_NEQ, 649), 	-- 516
is_word(IS_BRANCH, 648), 	-- 517
is_word(IS_READ, 249), 	-- 518
is_word(IS_SUB, 647), 	-- 519
is_word(IS_WRITE, 646), 	-- 520
is_word(IS_READ, 645), 	-- 521
is_word(IS_WRITE, 644), 	-- 522
is_word(IS_READ, 252), 	-- 523
is_word(IS_NEQ, 643), 	-- 524
is_word(IS_BRANCH, 642), 	-- 525
is_word(IS_READ, 249), 	-- 526
is_word(IS_ADD, 641), 	-- 527
is_word(IS_WRITE, 640), 	-- 528
is_word(IS_READ, 639), 	-- 529
is_word(IS_WRITE, 638), 	-- 530
is_word(IS_READ, 249), 	-- 531
is_word(IS_WRITE, 637), 	-- 532
is_word(IS_ADD, 3), 	-- 533
is_word(IS_WRITE, 636), 	-- 534
is_word(IS_READ, 635), 	-- 535
is_word(IS_WRITE, 2), 	-- 536
is_word(IS_READ, 249), 	-- 537
is_word(IS_WRITE, 2), 	-- 538
is_word(IS_READ, 634), 	-- 539
is_word(IS_WRITE, 2), 	-- 540
is_word(IS_READ, 633), 	-- 541
is_word(IS_WRITE, 632), 	-- 542
is_word(IS_READ, 2), 	-- 543
is_word(IS_WRITE, 631), 	-- 544
is_word(IS_ADD, 3), 	-- 545
is_word(IS_WRITE, 630), 	-- 546
is_word(IS_READ, 2), 	-- 547
is_word(IS_WRITE, 629), 	-- 548
is_word(IS_ADD, 3), 	-- 549
is_word(IS_WRITE, 628), 	-- 550
is_word(IS_READ, 253), 	-- 551
is_word(IS_EQ, 627), 	-- 552
is_word(IS_BRANCH, 626), 	-- 553
is_word(IS_READ, 253), 	-- 554
is_word(IS_SUB, 625), 	-- 555
is_word(IS_WRITE, 624), 	-- 556
is_word(IS_READ, 623), 	-- 557
is_word(IS_WRITE, 622), 	-- 558
is_word(IS_READ, 2), 	-- 559
is_word(IS_WRITE, 621), 	-- 560
is_word(IS_ADD, 3), 	-- 561
is_word(IS_WRITE, 620), 	-- 562
is_word(IS_READ, 2), 	-- 563
is_word(IS_WRITE, 619), 	-- 564
is_word(IS_ADD, 3), 	-- 565
is_word(IS_WRITE, 618), 	-- 566
is_word(IS_READ, 2), 	-- 567
is_word(IS_WRITE, 617), 	-- 568
is_word(IS_ADD, 3), 	-- 569
is_word(IS_WRITE, 616), 	-- 570
is_word(IS_READ, 254), 	-- 571
is_word(IS_WRITE, 615), 	-- 572
is_word(IS_ADD, 3), 	-- 573
is_word(IS_EQ, 614), 	-- 574
is_word(IS_BRANCH, 613), 	-- 575
is_word(IS_READ, 254), 	-- 576
is_word(IS_WRITE, 612), 	-- 577
is_word(IS_ADD, 3), 	-- 578
is_word(IS_WRITE, 255), 	-- 579
is_word(IS_READ, 254), 	-- 580
is_word(IS_ADD, 611), 	-- 581
is_word(IS_WRITE, 610), 	-- 582
is_word(IS_READ, 255), 	-- 583
is_word(IS_ADD, 609), 	-- 584
is_word(IS_WRITE, 608), 	-- 585
is_word(IS_READ, 607), 	-- 586
is_word(IS_WRITE, 606), 	-- 587
is_word(IS_READ, 2), 	-- 588
is_word(IS_WRITE, 605), 	-- 589
is_word(IS_ADD, 3), 	-- 590
is_word(IS_WRITE, 604), 	-- 591
0, 	-- 592
0, 	-- 593
0, 	-- 594
0, 	-- 595
0, 	-- 596
0, 	-- 597
0, 	-- 598
0, 	-- 599
0, 	-- 600
0, 	-- 601
0, 	-- 602
0, 	-- 603
0, 	-- 604
590, 	-- 605
0, 	-- 606
571, 	-- 607
255, 	-- 608
1, 	-- 609
254, 	-- 610
1, 	-- 611
578, 	-- 612
588, 	-- 613
0, 	-- 614
573, 	-- 615
255, 	-- 616
569, 	-- 617
254, 	-- 618
565, 	-- 619
0, 	-- 620
561, 	-- 621
0, 	-- 622
551, 	-- 623
253, 	-- 624
1, 	-- 625
559, 	-- 626
0, 	-- 627
253, 	-- 628
549, 	-- 629
0, 	-- 630
545, 	-- 631
0, 	-- 632
563, 	-- 633
337, 	-- 634
543, 	-- 635
248, 	-- 636
533, 	-- 637
0, 	-- 638
531, 	-- 639
249, 	-- 640
1, 	-- 641
531, 	-- 642
3, 	-- 643
0, 	-- 644
531, 	-- 645
249, 	-- 646
1, 	-- 647
523, 	-- 648
2, 	-- 649
0, 	-- 650
531, 	-- 651
249, 	-- 652
40, 	-- 653
515, 	-- 654
1, 	-- 655
0, 	-- 656
531, 	-- 657
249, 	-- 658
40, 	-- 659
507, 	-- 660
0, 	-- 661
249, 	-- 662
1104, 	-- 663
40, 	-- 664
252, 	-- 665
492, 	-- 666
251, 	-- 667
488, 	-- 668
250, 	-- 669
484, 	-- 670
0, 	-- 671
472, 	-- 672
1025, 	-- 673
48, 	-- 674
15, 	-- 675
1024, 	-- 676
48, 	-- 677
16, 	-- 678
0, 	-- 679
437, 	-- 680
196, 	-- 681
2, 	-- 682
0, 	-- 683
442, 	-- 684
197, 	-- 685
2, 	-- 686
445, 	-- 687
0, 	-- 688
482, 	-- 689
460, 	-- 690
445, 	-- 691
0, 	-- 692
192, 	-- 693
3, 	-- 694
467, 	-- 695
37, 	-- 696
197, 	-- 697
2, 	-- 698
472, 	-- 699
21, 	-- 700
196, 	-- 701
4, 	-- 702
0, 	-- 703
412, 	-- 704
196, 	-- 705
2, 	-- 706
415, 	-- 707
0, 	-- 708
482, 	-- 709
2, 	-- 710
428, 	-- 711
197, 	-- 712
3, 	-- 713
435, 	-- 714
37, 	-- 715
196, 	-- 716
2, 	-- 717
0, 	-- 718
360, 	-- 719
196, 	-- 720
1, 	-- 721
0, 	-- 722
365, 	-- 723
197, 	-- 724
1, 	-- 725
0, 	-- 726
563, 	-- 727
337, 	-- 728
400, 	-- 729
192, 	-- 730
1104, 	-- 731
40, 	-- 732
0, 	-- 733
400, 	-- 734
387, 	-- 735
0, 	-- 736
1, 	-- 737
387, 	-- 738
38, 	-- 739
387, 	-- 740
0, 	-- 741
387, 	-- 742
22, 	-- 743
387, 	-- 744
0, 	-- 745
405, 	-- 746
39, 	-- 747
197, 	-- 748
0, 	-- 749
410, 	-- 750
23, 	-- 751
196, 	-- 752
0, 	-- 753
355, 	-- 754
0, 	-- 755
0, 	-- 756
563, 	-- 757
326, 	-- 758
1104, 	-- 759
355, 	-- 760
0, 	-- 761
563, 	-- 762
290, 	-- 763
1024, 	-- 764
347, 	-- 765
0, 	-- 766
339	-- 767
